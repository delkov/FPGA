module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] addr,
    input go_home,
    // OUTPUT
    output [23:0] data,
    output rom_scan_is_done

  );
  
parameter rom_size = 4001;

reg [15:0] rom_data [rom_size:0];
reg [23:0] data_d, data_q;
wire[14:0] addrs;
reg [15:0] antidata;
reg done;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;


reg [15:0] CH_A_d, CH_A_q;
reg [15:0] CH_B_d, CH_B_q;
reg [15:0] CH_C_d, CH_C_q;
reg [15:0] CH_D_d, CH_D_q;


assign data = data_q;
assign rom_scan_is_done = done;
assign addrs = addr[15:2];


// always @(rst,addrs) begin
//   if (rst) begin
//       done = 1'b0;
//   end else begin
//       if (addrs == rom_size)
//           done = 1'b1;
//       else
//           done = 1'b0;
//   end     
// end // always
 

always @(*) begin
    
    CH_A_d=CH_A_q;
    CH_B_d=CH_B_q;
    CH_C_d=CH_C_q;
    CH_D_d=CH_D_q;

    if (go_home==1'b1) begin
        case (addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (CH_A_q>home_bias) begin
                    CH_A_d=CH_A_q-home_step;
                end else if (CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_A_d=CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (CH_C_q>home_bias) begin
                    CH_C_d=CH_C_q-home_step;
                end else if (CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_C_d=CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (CH_B_q>home_bias) begin
                    CH_B_d=CH_B_q-home_step;
                end else if (CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_B_d=CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (CH_D_q>home_bias) begin
                    CH_D_d=CH_D_q-home_step;
                end else if (CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_D_d=CH_D_q+home_step; 
                end 
            end

            default: begin
            end
        endcase

    end else begin // if go home==0
        case (addr[2:1])
            2'b00: begin
                CH_A_d= rom_data[addrs];
            end
            2'b01: begin
                CH_C_d= antidata;
            end
            2'b10: begin
                CH_B_d= rom_data[addrs];
            end
            2'b11: begin
                CH_D_d= antidata;
            end

        default: begin
            end
        endcase

    end // if go home 


    if (addrs == rom_size) begin
        done = 1'b1;
    end else begin
        done = 1'b0;
    end

end // always





always @(*) begin

    antidata = 16'hB900 - rom_data[addrs];
    
 
  rom_data[ 2]=16'b0010111101000111;
    rom_data[ 3]=16'b0101110111000000;
    rom_data[ 4]=16'b0010111101011100;
    rom_data[ 5]=16'b0101111100000100;
    rom_data[ 6]=16'b0010111101110001;
    rom_data[ 7]=16'b0110000001001000;
    rom_data[ 8]=16'b0010111110000110;
    rom_data[ 9]=16'b0110000110001100;
    rom_data[10]=16'b0010111110011011;
    rom_data[11]=16'b0110001011001111;
    rom_data[12]=16'b0010111110110000;
    rom_data[13]=16'b0110010000010010;
    rom_data[14]=16'b0010111111000101;
    rom_data[15]=16'b0110010101010100;
    rom_data[16]=16'b0010111111011010;
    rom_data[17]=16'b0110011010010101;
    rom_data[18]=16'b0010111111101111;
    rom_data[19]=16'b0110011111010101;
    rom_data[20]=16'b0011000000000100;
    rom_data[21]=16'b0110100100010101;
    rom_data[22]=16'b0011000000011010;
    rom_data[23]=16'b0110101001010011;
    rom_data[24]=16'b0011000000101111;
    rom_data[25]=16'b0110101110001111;
    rom_data[26]=16'b0011000001000101;
    rom_data[27]=16'b0110110011001011;
    rom_data[28]=16'b0011000001011011;
    rom_data[29]=16'b0110111000000100;
    rom_data[30]=16'b0011000001110001;
    rom_data[31]=16'b0110111100111100;
    rom_data[32]=16'b0011000010000111;
    rom_data[33]=16'b0111000001110010;
    rom_data[34]=16'b0011000010011101;
    rom_data[35]=16'b0111000110100110;
    rom_data[36]=16'b0011000010110011;
    rom_data[37]=16'b0111001011011000;
    rom_data[38]=16'b0011000011001010;
    rom_data[39]=16'b0111010000000111;
    rom_data[40]=16'b0011000011100001;
    rom_data[41]=16'b0111010100110011;
    rom_data[42]=16'b0011000011111000;
    rom_data[43]=16'b0111011001011101;
    rom_data[44]=16'b0011000100001111;
    rom_data[45]=16'b0111011110000011;
    rom_data[46]=16'b0011000100100110;
    rom_data[47]=16'b0111100010100110;
    rom_data[48]=16'b0011000100111110;
    rom_data[49]=16'b0111100111000110;
    rom_data[50]=16'b0011000101010110;
    rom_data[51]=16'b0111101011100001;
    rom_data[52]=16'b0011000101101110;
    rom_data[53]=16'b0111101111111001;
    rom_data[54]=16'b0011000110000111;
    rom_data[55]=16'b0111110100001011;
    rom_data[56]=16'b0011000110011111;
    rom_data[57]=16'b0111111000011001;
    rom_data[58]=16'b0011000110111000;
    rom_data[59]=16'b0111111100100010;
    rom_data[60]=16'b0011000111010001;
    rom_data[61]=16'b1000000000100101;
    rom_data[62]=16'b0011000111101011;
    rom_data[63]=16'b1000000100100010;
    rom_data[64]=16'b0011001000000101;
    rom_data[65]=16'b1000001000011001;
    rom_data[66]=16'b0011001000011111;
    rom_data[67]=16'b1000001100001001;
    rom_data[68]=16'b0011001000111010;
    rom_data[69]=16'b1000001111110010;
    rom_data[70]=16'b0011001001010100;
    rom_data[71]=16'b1000010011010010;
    rom_data[72]=16'b0011001001101111;
    rom_data[73]=16'b1000010110101010;
    rom_data[74]=16'b0011001010001011;
    rom_data[75]=16'b1000011001111001;
    rom_data[76]=16'b0011001010100111;
    rom_data[77]=16'b1000011100111110;
    rom_data[78]=16'b0011001011000010;
    rom_data[79]=16'b1000011111111001;
    rom_data[80]=16'b0011001011011111;
    rom_data[81]=16'b1000100010101001;
    rom_data[82]=16'b0011001011111011;
    rom_data[83]=16'b1000100101001110;
    rom_data[84]=16'b0011001100011000;
    rom_data[85]=16'b1000100111100101;
    rom_data[86]=16'b0011001100110101;
    rom_data[87]=16'b1000101001110000;
    rom_data[88]=16'b0011001101010010;
    rom_data[89]=16'b1000101011101101;
    rom_data[90]=16'b0011001101101111;
    rom_data[91]=16'b1000101101011011;
    rom_data[92]=16'b0011001110001100;
    rom_data[93]=16'b1000101110111010;
    rom_data[94]=16'b0011001110101001;
    rom_data[95]=16'b1000110000001010;
    rom_data[96]=16'b0011001111000110;
    rom_data[97]=16'b1000110001001001;
    rom_data[98]=16'b0011001111100100;
    rom_data[99]=16'b1000110001110111;
    rom_data[100]=16'b0011010000000001;
    rom_data[101]=16'b1000110010010100;
    rom_data[102]=16'b0011010000011101;
    rom_data[103]=16'b1000110010100000;
    rom_data[104]=16'b0011010000111010;
    rom_data[105]=16'b1000110010011010;
    rom_data[106]=16'b0011010001010111;
    rom_data[107]=16'b1000110010000011;
    rom_data[108]=16'b0011010001110011;
    rom_data[109]=16'b1000110001011010;
    rom_data[110]=16'b0011010010001111;
    rom_data[111]=16'b1000110000100001;
    rom_data[112]=16'b0011010010101011;
    rom_data[113]=16'b1000101111010110;
    rom_data[114]=16'b0011010011000110;
    rom_data[115]=16'b1000101101111011;
    rom_data[116]=16'b0011010011100001;
    rom_data[117]=16'b1000101100010001;
    rom_data[118]=16'b0011010011111100;
    rom_data[119]=16'b1000101010011000;
    rom_data[120]=16'b0011010100010111;
    rom_data[121]=16'b1000101000010000;
    rom_data[122]=16'b0011010100110001;
    rom_data[123]=16'b1000100101111010;
    rom_data[124]=16'b0011010101001011;
    rom_data[125]=16'b1000100011011000;
    rom_data[126]=16'b0011010101100101;
    rom_data[127]=16'b1000100000101001;
    rom_data[128]=16'b0011010101111110;
    rom_data[129]=16'b1000011101101110;
    rom_data[130]=16'b0011010110010111;
    rom_data[131]=16'b1000011010101001;
    rom_data[132]=16'b0011010110110000;
    rom_data[133]=16'b1000010111011010;
    rom_data[134]=16'b0011010111001000;
    rom_data[135]=16'b1000010100000001;
    rom_data[136]=16'b0011010111100001;
    rom_data[137]=16'b1000010000100000;
    rom_data[138]=16'b0011010111111000;
    rom_data[139]=16'b1000001100110110;
    rom_data[140]=16'b0011011000010000;
    rom_data[141]=16'b1000001001000101;
    rom_data[142]=16'b0011011000101000;
    rom_data[143]=16'b1000000101001101;
    rom_data[144]=16'b0011011000111111;
    rom_data[145]=16'b1000000001001110;
    rom_data[146]=16'b0011011001010110;
    rom_data[147]=16'b0111111101001001;
    rom_data[148]=16'b0011011001101101;
    rom_data[149]=16'b0111111000111110;
    rom_data[150]=16'b0011011010000011;
    rom_data[151]=16'b0111110100101110;
    rom_data[152]=16'b0011011010011010;
    rom_data[153]=16'b0111110000011001;
    rom_data[154]=16'b0011011010110000;
    rom_data[155]=16'b0111101100000000;
    rom_data[156]=16'b0011011011000110;
    rom_data[157]=16'b0111100111100010;
    rom_data[158]=16'b0011011011011100;
    rom_data[159]=16'b0111100011000000;
    rom_data[160]=16'b0011011011110010;
    rom_data[161]=16'b0111011110011011;
    rom_data[162]=16'b0011011100000111;
    rom_data[163]=16'b0111011001110011;
    rom_data[164]=16'b0011011100011101;
    rom_data[165]=16'b0111010101000111;
    rom_data[166]=16'b0011011100110010;
    rom_data[167]=16'b0111010000011001;
    rom_data[168]=16'b0011011101001000;
    rom_data[169]=16'b0111001011101000;
    rom_data[170]=16'b0011011101011101;
    rom_data[171]=16'b0111000110110101;
    rom_data[172]=16'b0011011101110010;
    rom_data[173]=16'b0111000001111111;
    rom_data[174]=16'b0011011110000111;
    rom_data[175]=16'b0110111101000111;
    rom_data[176]=16'b0011011110011100;
    rom_data[177]=16'b0110111000001110;
    rom_data[178]=16'b0011011110110001;
    rom_data[179]=16'b0110110011010011;
    rom_data[180]=16'b0011011111000110;
    rom_data[181]=16'b0110101110010110;
    rom_data[182]=16'b0011011111011011;
    rom_data[183]=16'b0110101001011000;
    rom_data[184]=16'b0011011111101111;
    rom_data[185]=16'b0110100100011001;
    rom_data[186]=16'b0011100000000100;
    rom_data[187]=16'b0110011111011001;
    rom_data[188]=16'b0011100000011001;
    rom_data[189]=16'b0110011010011000;
    rom_data[190]=16'b0011100000101101;
    rom_data[191]=16'b0110010101010110;
    rom_data[192]=16'b0011100001000010;
    rom_data[193]=16'b0110010000010011;
    rom_data[194]=16'b0011100001010111;
    rom_data[195]=16'b0110001011010000;
    rom_data[196]=16'b0011100001101011;
    rom_data[197]=16'b0110000110001100;
    rom_data[198]=16'b0011100010000000;
    rom_data[199]=16'b0110000001001000;
    rom_data[200]=16'b0011100010010101;
    rom_data[201]=16'b0101111100000100;
    rom_data[202]=16'b0011100010101001;
    rom_data[203]=16'b0101110111000000;
    rom_data[204]=16'b0011100010111110;
    rom_data[205]=16'b0101110001111100;
    rom_data[206]=16'b0011100011010011;
    rom_data[207]=16'b0101101100111000;
    rom_data[208]=16'b0011100011101000;
    rom_data[209]=16'b0101100111110100;
    rom_data[210]=16'b0011100011111101;
    rom_data[211]=16'b0101100010110001;
    rom_data[212]=16'b0011100100010010;
    rom_data[213]=16'b0101011101101110;
    rom_data[214]=16'b0011100100100111;
    rom_data[215]=16'b0101011000101100;
    rom_data[216]=16'b0011100100111100;
    rom_data[217]=16'b0101010011101011;
    rom_data[218]=16'b0011100101010001;
    rom_data[219]=16'b0101001110101011;
    rom_data[220]=16'b0011100101100110;
    rom_data[221]=16'b0101001001101011;
    rom_data[222]=16'b0011100101111100;
    rom_data[223]=16'b0101000100101101;
    rom_data[224]=16'b0011100110010001;
    rom_data[225]=16'b0100111111110000;
    rom_data[226]=16'b0011100110100111;
    rom_data[227]=16'b0100111010110101;
    rom_data[228]=16'b0011100110111101;
    rom_data[229]=16'b0100110101111011;
    rom_data[230]=16'b0011100111010011;
    rom_data[231]=16'b0100110001000011;
    rom_data[232]=16'b0011100111101001;
    rom_data[233]=16'b0100101100001101;
    rom_data[234]=16'b0011100111111111;
    rom_data[235]=16'b0100100111011010;
    rom_data[236]=16'b0011101000010101;
    rom_data[237]=16'b0100100010101000;
    rom_data[238]=16'b0011101000101100;
    rom_data[239]=16'b0100011101111001;
    rom_data[240]=16'b0011101001000011;
    rom_data[241]=16'b0100011001001100;
    rom_data[242]=16'b0011101001011010;
    rom_data[243]=16'b0100010100100011;
    rom_data[244]=16'b0011101001110001;
    rom_data[245]=16'b0100001111111100;
    rom_data[246]=16'b0011101010001000;
    rom_data[247]=16'b0100001011011001;
    rom_data[248]=16'b0011101010100000;
    rom_data[249]=16'b0100000110111010;
    rom_data[250]=16'b0011101010111000;
    rom_data[251]=16'b0100000010011111;
    rom_data[252]=16'b0011101011010000;
    rom_data[253]=16'b0011111110000111;
    rom_data[254]=16'b0011101011101001;
    rom_data[255]=16'b0011111001110100;
    rom_data[256]=16'b0011101100000001;
    rom_data[257]=16'b0011110101100110;
    rom_data[258]=16'b0011101100011010;
    rom_data[259]=16'b0011110001011110;
    rom_data[260]=16'b0011101100110100;
    rom_data[261]=16'b0011101101011011;
    rom_data[262]=16'b0011101101001101;
    rom_data[263]=16'b0011101001011101;
    rom_data[264]=16'b0011101101100111;
    rom_data[265]=16'b0011100101100111;
    rom_data[266]=16'b0011101110000001;
    rom_data[267]=16'b0011100001110111;
    rom_data[268]=16'b0011101110011100;
    rom_data[269]=16'b0011011110001110;
    rom_data[270]=16'b0011101110110110;
    rom_data[271]=16'b0011011010101110;
    rom_data[272]=16'b0011101111010010;
    rom_data[273]=16'b0011010111010110;
    rom_data[274]=16'b0011101111101101;
    rom_data[275]=16'b0011010100000111;
    rom_data[276]=16'b0011110000001001;
    rom_data[277]=16'b0011010001000001;
    rom_data[278]=16'b0011110000100101;
    rom_data[279]=16'b0011001110000111;
    rom_data[280]=16'b0011110001000001;
    rom_data[281]=16'b0011001011010111;
    rom_data[282]=16'b0011110001011101;
    rom_data[283]=16'b0011001000110010;
    rom_data[284]=16'b0011110001111010;
    rom_data[285]=16'b0011000110011011;
    rom_data[286]=16'b0011110010010111;
    rom_data[287]=16'b0011000100010000;
    rom_data[288]=16'b0011110010110100;
    rom_data[289]=16'b0011000010010011;
    rom_data[290]=16'b0011110011010001;
    rom_data[291]=16'b0011000000100101;
    rom_data[292]=16'b0011110011101110;
    rom_data[293]=16'b0010111111000110;
    rom_data[294]=16'b0011110100001011;
    rom_data[295]=16'b0010111101110110;
    rom_data[296]=16'b0011110100101000;
    rom_data[297]=16'b0010111100110111;
    rom_data[298]=16'b0011110101000110;
    rom_data[299]=16'b0010111100001001;
    rom_data[300]=16'b0011110101100011;
    rom_data[301]=16'b0010111011101100;
    rom_data[302]=16'b0011110110000000;
    rom_data[303]=16'b0010111011100000;
    rom_data[304]=16'b0011110110011100;
    rom_data[305]=16'b0010111011100110;
    rom_data[306]=16'b0011110110111001;
    rom_data[307]=16'b0010111011111101;
    rom_data[308]=16'b0011110111010101;
    rom_data[309]=16'b0010111100100110;
    rom_data[310]=16'b0011110111110001;
    rom_data[311]=16'b0010111101011111;
    rom_data[312]=16'b0011111000001101;
    rom_data[313]=16'b0010111110101010;
    rom_data[314]=16'b0011111000101000;
    rom_data[315]=16'b0011000000000101;
    rom_data[316]=16'b0011111001000100;
    rom_data[317]=16'b0011000001101111;
    rom_data[318]=16'b0011111001011110;
    rom_data[319]=16'b0011000011101000;
    rom_data[320]=16'b0011111001111001;
    rom_data[321]=16'b0011000101110000;
    rom_data[322]=16'b0011111010010011;
    rom_data[323]=16'b0011001000000110;
    rom_data[324]=16'b0011111010101101;
    rom_data[325]=16'b0011001010101001;
    rom_data[326]=16'b0011111011000111;
    rom_data[327]=16'b0011001101010111;
    rom_data[328]=16'b0011111011100000;
    rom_data[329]=16'b0011010000010010;
    rom_data[330]=16'b0011111011111001;
    rom_data[331]=16'b0011010011010111;
    rom_data[332]=16'b0011111100010010;
    rom_data[333]=16'b0011010110100110;
    rom_data[334]=16'b0011111100101010;
    rom_data[335]=16'b0011011001111111;
    rom_data[336]=16'b0011111101000011;
    rom_data[337]=16'b0011011101100000;
    rom_data[338]=16'b0011111101011011;
    rom_data[339]=16'b0011100001001010;
    rom_data[340]=16'b0011111101110010;
    rom_data[341]=16'b0011100100111011;
    rom_data[342]=16'b0011111110001010;
    rom_data[343]=16'b0011101000110100;
    rom_data[344]=16'b0011111110100001;
    rom_data[345]=16'b0011101100110010;
    rom_data[346]=16'b0011111110111000;
    rom_data[347]=16'b0011110000111000;
    rom_data[348]=16'b0011111111001111;
    rom_data[349]=16'b0011110101000010;
    rom_data[350]=16'b0011111111100101;
    rom_data[351]=16'b0011111001010010;
    rom_data[352]=16'b0011111111111100;
    rom_data[353]=16'b0011111101100111;
    rom_data[354]=16'b0100000000010010;
    rom_data[355]=16'b0100000010000001;
    rom_data[356]=16'b0100000000101000;
    rom_data[357]=16'b0100000110011110;
    rom_data[358]=16'b0100000000111110;
    rom_data[359]=16'b0100001011000000;
    rom_data[360]=16'b0100000001010100;
    rom_data[361]=16'b0100001111100101;
    rom_data[362]=16'b0100000001101010;
    rom_data[363]=16'b0100010100001101;
    rom_data[364]=16'b0100000001111111;
    rom_data[365]=16'b0100011000111001;
    rom_data[366]=16'b0100000010010100;
    rom_data[367]=16'b0100011101100111;
    rom_data[368]=16'b0100000010101010;
    rom_data[369]=16'b0100100010011000;
    rom_data[370]=16'b0100000010111111;
    rom_data[371]=16'b0100100111001011;
    rom_data[372]=16'b0100000011010100;
    rom_data[373]=16'b0100101100000001;
    rom_data[374]=16'b0100000011101001;
    rom_data[375]=16'b0100110000111001;
    rom_data[376]=16'b0100000011111110;
    rom_data[377]=16'b0100110101110010;
    rom_data[378]=16'b0100000100010011;
    rom_data[379]=16'b0100111010101101;
    rom_data[380]=16'b0100000100101000;
    rom_data[381]=16'b0100111111101010;
    rom_data[382]=16'b0100000100111101;
    rom_data[383]=16'b0101000100101000;
    rom_data[384]=16'b0100000101010001;
    rom_data[385]=16'b0101001001100111;
    rom_data[386]=16'b0100000101100110;
    rom_data[387]=16'b0101001110100111;
    rom_data[388]=16'b0100000101111011;
    rom_data[389]=16'b0101010011101001;
    rom_data[390]=16'b0100000110001111;
    rom_data[391]=16'b0101011000101011;
    rom_data[392]=16'b0100000110100100;
    rom_data[393]=16'b0101011101101101;
    rom_data[394]=16'b0100000110111001;
    rom_data[395]=16'b0101100010110001;
    rom_data[396]=16'b0100000111001101;
    rom_data[397]=16'b0101100111110100;
    rom_data[398]=16'b0100000111100010;
    rom_data[399]=16'b0101101100111000;
    rom_data[400]=16'b0100000111110111;
    rom_data[401]=16'b0101110001111100;
    rom_data[402]=16'b0100001000001100;
    rom_data[403]=16'b0101110111000000;
    rom_data[404]=16'b0100001000100000;
    rom_data[405]=16'b0101111100000100;
    rom_data[406]=16'b0100001000110101;
    rom_data[407]=16'b0110000001001000;
    rom_data[408]=16'b0100001001001010;
    rom_data[409]=16'b0110000110001100;
    rom_data[410]=16'b0100001001011111;
    rom_data[411]=16'b0110001011001111;
    rom_data[412]=16'b0100001001110100;
    rom_data[413]=16'b0110010000010010;
    rom_data[414]=16'b0100001010001001;
    rom_data[415]=16'b0110010101010100;
    rom_data[416]=16'b0100001010011110;
    rom_data[417]=16'b0110011010010101;
    rom_data[418]=16'b0100001010110011;
    rom_data[419]=16'b0110011111010110;
    rom_data[420]=16'b0100001011001000;
    rom_data[421]=16'b0110100100010101;
    rom_data[422]=16'b0100001011011110;
    rom_data[423]=16'b0110101001010011;
    rom_data[424]=16'b0100001011110011;
    rom_data[425]=16'b0110101110010000;
    rom_data[426]=16'b0100001100001001;
    rom_data[427]=16'b0110110011001011;
    rom_data[428]=16'b0100001100011111;
    rom_data[429]=16'b0110111000000101;
    rom_data[430]=16'b0100001100110101;
    rom_data[431]=16'b0110111100111101;
    rom_data[432]=16'b0100001101001011;
    rom_data[433]=16'b0111000001110011;
    rom_data[434]=16'b0100001101100001;
    rom_data[435]=16'b0111000110100111;
    rom_data[436]=16'b0100001101110111;
    rom_data[437]=16'b0111001011011000;
    rom_data[438]=16'b0100001110001110;
    rom_data[439]=16'b0111010000000111;
    rom_data[440]=16'b0100001110100101;
    rom_data[441]=16'b0111010100110100;
    rom_data[442]=16'b0100001110111100;
    rom_data[443]=16'b0111011001011101;
    rom_data[444]=16'b0100001111010011;
    rom_data[445]=16'b0111011110000100;
    rom_data[446]=16'b0100001111101010;
    rom_data[447]=16'b0111100010100111;
    rom_data[448]=16'b0100010000000010;
    rom_data[449]=16'b0111100111000110;
    rom_data[450]=16'b0100010000011010;
    rom_data[451]=16'b0111101011100010;
    rom_data[452]=16'b0100010000110010;
    rom_data[453]=16'b0111101111111001;
    rom_data[454]=16'b0100010001001011;
    rom_data[455]=16'b0111110100001100;
    rom_data[456]=16'b0100010001100011;
    rom_data[457]=16'b0111111000011010;
    rom_data[458]=16'b0100010001111100;
    rom_data[459]=16'b0111111100100010;
    rom_data[460]=16'b0100010010010110;
    rom_data[461]=16'b1000000000100110;
    rom_data[462]=16'b0100010010101111;
    rom_data[463]=16'b1000000100100011;
    rom_data[464]=16'b0100010011001001;
    rom_data[465]=16'b1000001000011010;
    rom_data[466]=16'b0100010011100011;
    rom_data[467]=16'b1000001100001001;
    rom_data[468]=16'b0100010011111110;
    rom_data[469]=16'b1000001111110010;
    rom_data[470]=16'b0100010100011000;
    rom_data[471]=16'b1000010011010010;
    rom_data[472]=16'b0100010100110100;
    rom_data[473]=16'b1000010110101010;
    rom_data[474]=16'b0100010101001111;
    rom_data[475]=16'b1000011001111001;
    rom_data[476]=16'b0100010101101011;
    rom_data[477]=16'b1000011100111111;
    rom_data[478]=16'b0100010110000111;
    rom_data[479]=16'b1000011111111010;
    rom_data[480]=16'b0100010110100011;
    rom_data[481]=16'b1000100010101010;
    rom_data[482]=16'b0100010110111111;
    rom_data[483]=16'b1000100101001110;
    rom_data[484]=16'b0100010111011100;
    rom_data[485]=16'b1000100111100110;
    rom_data[486]=16'b0100010111111001;
    rom_data[487]=16'b1000101001110000;
    rom_data[488]=16'b0100011000010110;
    rom_data[489]=16'b1000101011101101;
    rom_data[490]=16'b0100011000110011;
    rom_data[491]=16'b1000101101011011;
    rom_data[492]=16'b0100011001010000;
    rom_data[493]=16'b1000101110111010;
    rom_data[494]=16'b0100011001101101;
    rom_data[495]=16'b1000110000001010;
    rom_data[496]=16'b0100011010001011;
    rom_data[497]=16'b1000110001001001;
    rom_data[498]=16'b0100011010101000;
    rom_data[499]=16'b1000110001110111;
    rom_data[500]=16'b0100011011000101;
    rom_data[501]=16'b1000110010010100;
    rom_data[502]=16'b0100011011100010;
    rom_data[503]=16'b1000110010100000;
    rom_data[504]=16'b0100011011111110;
    rom_data[505]=16'b1000110010011010;
    rom_data[506]=16'b0100011100011011;
    rom_data[507]=16'b1000110010000011;
    rom_data[508]=16'b0100011100110111;
    rom_data[509]=16'b1000110001011010;
    rom_data[510]=16'b0100011101010011;
    rom_data[511]=16'b1000110000100000;
    rom_data[512]=16'b0100011101101111;
    rom_data[513]=16'b1000101111010110;
    rom_data[514]=16'b0100011110001010;
    rom_data[515]=16'b1000101101111011;
    rom_data[516]=16'b0100011110100110;
    rom_data[517]=16'b1000101100010001;
    rom_data[518]=16'b0100011111000001;
    rom_data[519]=16'b1000101010010111;
    rom_data[520]=16'b0100011111011011;
    rom_data[521]=16'b1000101000010000;
    rom_data[522]=16'b0100011111110101;
    rom_data[523]=16'b1000100101111010;
    rom_data[524]=16'b0100100000001111;
    rom_data[525]=16'b1000100011010111;
    rom_data[526]=16'b0100100000101001;
    rom_data[527]=16'b1000100000101000;
    rom_data[528]=16'b0100100001000010;
    rom_data[529]=16'b1000011101101110;
    rom_data[530]=16'b0100100001011011;
    rom_data[531]=16'b1000011010101001;
    rom_data[532]=16'b0100100001110100;
    rom_data[533]=16'b1000010111011010;
    rom_data[534]=16'b0100100010001100;
    rom_data[535]=16'b1000010100000001;
    rom_data[536]=16'b0100100010100101;
    rom_data[537]=16'b1000010000100000;
    rom_data[538]=16'b0100100010111101;
    rom_data[539]=16'b1000001100110110;
    rom_data[540]=16'b0100100011010100;
    rom_data[541]=16'b1000001001000101;
    rom_data[542]=16'b0100100011101100;
    rom_data[543]=16'b1000000101001100;
    rom_data[544]=16'b0100100100000011;
    rom_data[545]=16'b1000000001001101;
    rom_data[546]=16'b0100100100011010;
    rom_data[547]=16'b0111111101001000;
    rom_data[548]=16'b0100100100110001;
    rom_data[549]=16'b0111111000111110;
    rom_data[550]=16'b0100100101000111;
    rom_data[551]=16'b0111110100101110;
    rom_data[552]=16'b0100100101011110;
    rom_data[553]=16'b0111110000011001;
    rom_data[554]=16'b0100100101110100;
    rom_data[555]=16'b0111101011111111;
    rom_data[556]=16'b0100100110001010;
    rom_data[557]=16'b0111100111100010;
    rom_data[558]=16'b0100100110100000;
    rom_data[559]=16'b0111100011000000;
    rom_data[560]=16'b0100100110110110;
    rom_data[561]=16'b0111011110011011;
    rom_data[562]=16'b0100100111001100;
    rom_data[563]=16'b0111011001110011;
    rom_data[564]=16'b0100100111100001;
    rom_data[565]=16'b0111010101000111;
    rom_data[566]=16'b0100100111110111;
    rom_data[567]=16'b0111010000011001;
    rom_data[568]=16'b0100101000001100;
    rom_data[569]=16'b0111001011101000;
    rom_data[570]=16'b0100101000100001;
    rom_data[571]=16'b0111000110110100;
    rom_data[572]=16'b0100101000110110;
    rom_data[573]=16'b0111000001111111;
    rom_data[574]=16'b0100101001001011;
    rom_data[575]=16'b0110111101000111;
    rom_data[576]=16'b0100101001100000;
    rom_data[577]=16'b0110111000001110;
    rom_data[578]=16'b0100101001110101;
    rom_data[579]=16'b0110110011010011;
    rom_data[580]=16'b0100101010001010;
    rom_data[581]=16'b0110101110010110;
    rom_data[582]=16'b0100101010011111;
    rom_data[583]=16'b0110101001011000;
    rom_data[584]=16'b0100101010110011;
    rom_data[585]=16'b0110100100011001;
    rom_data[586]=16'b0100101011001000;
    rom_data[587]=16'b0110011111011000;
    rom_data[588]=16'b0100101011011101;
    rom_data[589]=16'b0110011010010111;
    rom_data[590]=16'b0100101011110010;
    rom_data[591]=16'b0110010101010101;
    rom_data[592]=16'b0100101100000110;
    rom_data[593]=16'b0110010000010011;
    rom_data[594]=16'b0100101100011011;
    rom_data[595]=16'b0110001011001111;
    rom_data[596]=16'b0100101100110000;
    rom_data[597]=16'b0110000110001100;
    rom_data[598]=16'b0100101101000100;
    rom_data[599]=16'b0110000001001000;
    rom_data[600]=16'b0100101101011001;
    rom_data[601]=16'b0101111100000100;
    rom_data[602]=16'b0100101101101110;
    rom_data[603]=16'b0101110110111111;
    rom_data[604]=16'b0100101110000010;
    rom_data[605]=16'b0101110001111011;
    rom_data[606]=16'b0100101110010111;
    rom_data[607]=16'b0101101100110111;
    rom_data[608]=16'b0100101110101100;
    rom_data[609]=16'b0101100111110100;
    rom_data[610]=16'b0100101111000001;
    rom_data[611]=16'b0101100010110001;
    rom_data[612]=16'b0100101111010110;
    rom_data[613]=16'b0101011101101110;
    rom_data[614]=16'b0100101111101011;
    rom_data[615]=16'b0101011000101100;
    rom_data[616]=16'b0100110000000000;
    rom_data[617]=16'b0101010011101011;
    rom_data[618]=16'b0100110000010101;
    rom_data[619]=16'b0101001110101010;
    rom_data[620]=16'b0100110000101010;
    rom_data[621]=16'b0101001001101011;
    rom_data[622]=16'b0100110001000000;
    rom_data[623]=16'b0101000100101101;
    rom_data[624]=16'b0100110001010101;
    rom_data[625]=16'b0100111111110000;
    rom_data[626]=16'b0100110001101011;
    rom_data[627]=16'b0100111010110101;
    rom_data[628]=16'b0100110010000001;
    rom_data[629]=16'b0100110101111011;
    rom_data[630]=16'b0100110010010111;
    rom_data[631]=16'b0100110001000011;
    rom_data[632]=16'b0100110010101101;
    rom_data[633]=16'b0100101100001101;
    rom_data[634]=16'b0100110011000011;
    rom_data[635]=16'b0100100111011001;
    rom_data[636]=16'b0100110011011010;
    rom_data[637]=16'b0100100010101000;
    rom_data[638]=16'b0100110011110000;
    rom_data[639]=16'b0100011101111000;
    rom_data[640]=16'b0100110100000111;
    rom_data[641]=16'b0100011001001100;
    rom_data[642]=16'b0100110100011110;
    rom_data[643]=16'b0100010100100011;
    rom_data[644]=16'b0100110100110101;
    rom_data[645]=16'b0100001111111100;
    rom_data[646]=16'b0100110101001101;
    rom_data[647]=16'b0100001011011001;
    rom_data[648]=16'b0100110101100100;
    rom_data[649]=16'b0100000110111010;
    rom_data[650]=16'b0100110101111100;
    rom_data[651]=16'b0100000010011110;
    rom_data[652]=16'b0100110110010100;
    rom_data[653]=16'b0011111110000111;
    rom_data[654]=16'b0100110110101101;
    rom_data[655]=16'b0011111001110100;
    rom_data[656]=16'b0100110111000101;
    rom_data[657]=16'b0011110101100110;
    rom_data[658]=16'b0100110111011110;
    rom_data[659]=16'b0011110001011101;
    rom_data[660]=16'b0100110111111000;
    rom_data[661]=16'b0011101101011010;
    rom_data[662]=16'b0100111000010001;
    rom_data[663]=16'b0011101001011101;
    rom_data[664]=16'b0100111000101011;
    rom_data[665]=16'b0011100101100110;
    rom_data[666]=16'b0100111001000101;
    rom_data[667]=16'b0011100001110111;
    rom_data[668]=16'b0100111001100000;
    rom_data[669]=16'b0011011110001110;
    rom_data[670]=16'b0100111001111011;
    rom_data[671]=16'b0011011010101110;
    rom_data[672]=16'b0100111010010110;
    rom_data[673]=16'b0011010111010101;
    rom_data[674]=16'b0100111010110001;
    rom_data[675]=16'b0011010100000111;
    rom_data[676]=16'b0100111011001101;
    rom_data[677]=16'b0011010001000001;
    rom_data[678]=16'b0100111011101001;
    rom_data[679]=16'b0011001110000110;
    rom_data[680]=16'b0100111100000101;
    rom_data[681]=16'b0011001011010110;
    rom_data[682]=16'b0100111100100001;
    rom_data[683]=16'b0011001000110010;
    rom_data[684]=16'b0100111100111110;
    rom_data[685]=16'b0011000110011010;
    rom_data[686]=16'b0100111101011011;
    rom_data[687]=16'b0011000100010000;
    rom_data[688]=16'b0100111101111000;
    rom_data[689]=16'b0011000010010011;
    rom_data[690]=16'b0100111110010101;
    rom_data[691]=16'b0011000000100101;
    rom_data[692]=16'b0100111110110010;
    rom_data[693]=16'b0010111111000110;
    rom_data[694]=16'b0100111111001111;
    rom_data[695]=16'b0010111101110110;
    rom_data[696]=16'b0100111111101101;
    rom_data[697]=16'b0010111100110111;
    rom_data[698]=16'b0101000000001010;
    rom_data[699]=16'b0010111100001001;
    rom_data[700]=16'b0101000000100111;
    rom_data[701]=16'b0010111011101100;
    rom_data[702]=16'b0101000001000100;
    rom_data[703]=16'b0010111011100000;
    rom_data[704]=16'b0101000001100000;
    rom_data[705]=16'b0010111011100110;
    rom_data[706]=16'b0101000001111101;
    rom_data[707]=16'b0010111011111101;
    rom_data[708]=16'b0101000010011001;
    rom_data[709]=16'b0010111100100110;
    rom_data[710]=16'b0101000010110101;
    rom_data[711]=16'b0010111101100000;
    rom_data[712]=16'b0101000011010001;
    rom_data[713]=16'b0010111110101010;
    rom_data[714]=16'b0101000011101101;
    rom_data[715]=16'b0011000000000101;
    rom_data[716]=16'b0101000100001000;
    rom_data[717]=16'b0011000001101111;
    rom_data[718]=16'b0101000100100011;
    rom_data[719]=16'b0011000011101001;
    rom_data[720]=16'b0101000100111101;
    rom_data[721]=16'b0011000101110001;
    rom_data[722]=16'b0101000101010111;
    rom_data[723]=16'b0011001000000110;
    rom_data[724]=16'b0101000101110001;
    rom_data[725]=16'b0011001010101001;
    rom_data[726]=16'b0101000110001011;
    rom_data[727]=16'b0011001101011000;
    rom_data[728]=16'b0101000110100100;
    rom_data[729]=16'b0011010000010010;
    rom_data[730]=16'b0101000110111101;
    rom_data[731]=16'b0011010011010111;
    rom_data[732]=16'b0101000111010110;
    rom_data[733]=16'b0011010110100110;
    rom_data[734]=16'b0101000111101111;
    rom_data[735]=16'b0011011001111111;
    rom_data[736]=16'b0101001000000111;
    rom_data[737]=16'b0011011101100000;
    rom_data[738]=16'b0101001000011111;
    rom_data[739]=16'b0011100001001010;
    rom_data[740]=16'b0101001000110110;
    rom_data[741]=16'b0011100100111011;
    rom_data[742]=16'b0101001001001110;
    rom_data[743]=16'b0011101000110100;
    rom_data[744]=16'b0101001001100101;
    rom_data[745]=16'b0011101100110011;
    rom_data[746]=16'b0101001001111100;
    rom_data[747]=16'b0011110000111000;
    rom_data[748]=16'b0101001010010011;
    rom_data[749]=16'b0011110101000011;
    rom_data[750]=16'b0101001010101010;
    rom_data[751]=16'b0011111001010011;
    rom_data[752]=16'b0101001011000000;
    rom_data[753]=16'b0011111101100111;
    rom_data[754]=16'b0101001011010110;
    rom_data[755]=16'b0100000010000001;
    rom_data[756]=16'b0101001011101100;
    rom_data[757]=16'b0100000110011111;
    rom_data[758]=16'b0101001100000010;
    rom_data[759]=16'b0100001011000000;
    rom_data[760]=16'b0101001100011000;
    rom_data[761]=16'b0100001111100101;
    rom_data[762]=16'b0101001100101110;
    rom_data[763]=16'b0100010100001110;
    rom_data[764]=16'b0101001101000011;
    rom_data[765]=16'b0100011000111001;
    rom_data[766]=16'b0101001101011001;
    rom_data[767]=16'b0100011101100111;
    rom_data[768]=16'b0101001101101110;
    rom_data[769]=16'b0100100010011000;
    rom_data[770]=16'b0101001110000011;
    rom_data[771]=16'b0100100111001100;
    rom_data[772]=16'b0101001110011000;
    rom_data[773]=16'b0100101100000001;
    rom_data[774]=16'b0101001110101101;
    rom_data[775]=16'b0100110000111001;
    rom_data[776]=16'b0101001111000010;
    rom_data[777]=16'b0100110101110011;
    rom_data[778]=16'b0101001111010111;
    rom_data[779]=16'b0100111010101110;
    rom_data[780]=16'b0101001111101100;
    rom_data[781]=16'b0100111111101010;
    rom_data[782]=16'b0101010000000001;
    rom_data[783]=16'b0101000100101000;
    rom_data[784]=16'b0101010000010110;
    rom_data[785]=16'b0101001001100111;
    rom_data[786]=16'b0101010000101010;
    rom_data[787]=16'b0101001110101000;
    rom_data[788]=16'b0101010000111111;
    rom_data[789]=16'b0101010011101001;
    rom_data[790]=16'b0101010001010100;
    rom_data[791]=16'b0101011000101011;
    rom_data[792]=16'b0101010001101000;
    rom_data[793]=16'b0101011101101110;
    rom_data[794]=16'b0101010001111101;
    rom_data[795]=16'b0101100010110001;
    rom_data[796]=16'b0101010010010010;
    rom_data[797]=16'b0101100111110101;
    rom_data[798]=16'b0101010010100110;
    rom_data[799]=16'b0101101100111000;
    rom_data[800]=16'b0101010010111011;
    rom_data[801]=16'b0101110001111101;
    rom_data[802]=16'b0101010011010000;
    rom_data[803]=16'b0101110111000001;
    rom_data[804]=16'b0101010011100100;
    rom_data[805]=16'b0101111100000101;
    rom_data[806]=16'b0101010011111001;
    rom_data[807]=16'b0110000001001001;
    rom_data[808]=16'b0101010100001110;
    rom_data[809]=16'b0110000110001100;
    rom_data[810]=16'b0101010100100011;
    rom_data[811]=16'b0110001011010000;
    rom_data[812]=16'b0101010100111000;
    rom_data[813]=16'b0110010000010010;
    rom_data[814]=16'b0101010101001101;
    rom_data[815]=16'b0110010101010100;
    rom_data[816]=16'b0101010101100010;
    rom_data[817]=16'b0110011010010110;
    rom_data[818]=16'b0101010101110111;
    rom_data[819]=16'b0110011111010110;
    rom_data[820]=16'b0101010110001101;
    rom_data[821]=16'b0110100100010101;
    rom_data[822]=16'b0101010110100010;
    rom_data[823]=16'b0110101001010011;
    rom_data[824]=16'b0101010110110111;
    rom_data[825]=16'b0110101110010000;
    rom_data[826]=16'b0101010111001101;
    rom_data[827]=16'b0110110011001011;
    rom_data[828]=16'b0101010111100011;
    rom_data[829]=16'b0110111000000101;
    rom_data[830]=16'b0101010111111001;
    rom_data[831]=16'b0110111100111101;
    rom_data[832]=16'b0101011000001111;
    rom_data[833]=16'b0111000001110011;
    rom_data[834]=16'b0101011000100101;
    rom_data[835]=16'b0111000110100111;
    rom_data[836]=16'b0101011000111100;
    rom_data[837]=16'b0111001011011001;
    rom_data[838]=16'b0101011001010010;
    rom_data[839]=16'b0111010000001000;
    rom_data[840]=16'b0101011001101001;
    rom_data[841]=16'b0111010100110100;
    rom_data[842]=16'b0101011010000000;
    rom_data[843]=16'b0111011001011110;
    rom_data[844]=16'b0101011010010111;
    rom_data[845]=16'b0111011110000100;
    rom_data[846]=16'b0101011010101111;
    rom_data[847]=16'b0111100010100111;
    rom_data[848]=16'b0101011011000110;
    rom_data[849]=16'b0111100111000110;
    rom_data[850]=16'b0101011011011110;
    rom_data[851]=16'b0111101011100010;
    rom_data[852]=16'b0101011011110110;
    rom_data[853]=16'b0111101111111001;
    rom_data[854]=16'b0101011100001111;
    rom_data[855]=16'b0111110100001100;
    rom_data[856]=16'b0101011100100111;
    rom_data[857]=16'b0111111000011010;
    rom_data[858]=16'b0101011101000000;
    rom_data[859]=16'b0111111100100011;
    rom_data[860]=16'b0101011101011010;
    rom_data[861]=16'b1000000000100110;
    rom_data[862]=16'b0101011101110011;
    rom_data[863]=16'b1000000100100011;
    rom_data[864]=16'b0101011110001101;
    rom_data[865]=16'b1000001000011010;
    rom_data[866]=16'b0101011110100111;
    rom_data[867]=16'b1000001100001010;
    rom_data[868]=16'b0101011111000010;
    rom_data[869]=16'b1000001111110010;
    rom_data[870]=16'b0101011111011101;
    rom_data[871]=16'b1000010011010011;
    rom_data[872]=16'b0101011111111000;
    rom_data[873]=16'b1000010110101011;
    rom_data[874]=16'b0101100000010011;
    rom_data[875]=16'b1000011001111010;
    rom_data[876]=16'b0101100000101111;
    rom_data[877]=16'b1000011100111111;
    rom_data[878]=16'b0101100001001011;
    rom_data[879]=16'b1000011111111010;
    rom_data[880]=16'b0101100001100111;
    rom_data[881]=16'b1000100010101010;
    rom_data[882]=16'b0101100010000011;
    rom_data[883]=16'b1000100101001110;
    rom_data[884]=16'b0101100010100000;
    rom_data[885]=16'b1000100111100110;
    rom_data[886]=16'b0101100010111101;
    rom_data[887]=16'b1000101001110000;
    rom_data[888]=16'b0101100011011010;
    rom_data[889]=16'b1000101011101101;
    rom_data[890]=16'b0101100011110111;
    rom_data[891]=16'b1000101101011011;
    rom_data[892]=16'b0101100100010100;
    rom_data[893]=16'b1000101110111010;
    rom_data[894]=16'b0101100100110001;
    rom_data[895]=16'b1000110000001010;
    rom_data[896]=16'b0101100101001111;
    rom_data[897]=16'b1000110001001001;
    rom_data[898]=16'b0101100101101100;
    rom_data[899]=16'b1000110001110111;
    rom_data[900]=16'b0101100110001001;
    rom_data[901]=16'b1000110010010100;
    rom_data[902]=16'b0101100110100110;
    rom_data[903]=16'b1000110010100000;
    rom_data[904]=16'b0101100111000010;
    rom_data[905]=16'b1000110010011010;
    rom_data[906]=16'b0101100111011111;
    rom_data[907]=16'b1000110010000011;
    rom_data[908]=16'b0101100111111011;
    rom_data[909]=16'b1000110001011010;
    rom_data[910]=16'b0101101000010111;
    rom_data[911]=16'b1000110000100000;
    rom_data[912]=16'b0101101000110011;
    rom_data[913]=16'b1000101111010110;
    rom_data[914]=16'b0101101001001111;
    rom_data[915]=16'b1000101101111011;
    rom_data[916]=16'b0101101001101010;
    rom_data[917]=16'b1000101100010001;
    rom_data[918]=16'b0101101010000101;
    rom_data[919]=16'b1000101010010111;
    rom_data[920]=16'b0101101010011111;
    rom_data[921]=16'b1000101000001111;
    rom_data[922]=16'b0101101010111001;
    rom_data[923]=16'b1000100101111010;
    rom_data[924]=16'b0101101011010011;
    rom_data[925]=16'b1000100011010111;
    rom_data[926]=16'b0101101011101101;
    rom_data[927]=16'b1000100000101000;
    rom_data[928]=16'b0101101100000110;
    rom_data[929]=16'b1000011101101110;
    rom_data[930]=16'b0101101100011111;
    rom_data[931]=16'b1000011010101001;
    rom_data[932]=16'b0101101100111000;
    rom_data[933]=16'b1000010111011010;
    rom_data[934]=16'b0101101101010001;
    rom_data[935]=16'b1000010100000001;
    rom_data[936]=16'b0101101101101001;
    rom_data[937]=16'b1000010000011111;
    rom_data[938]=16'b0101101110000001;
    rom_data[939]=16'b1000001100110110;
    rom_data[940]=16'b0101101110011000;
    rom_data[941]=16'b1000001001000100;
    rom_data[942]=16'b0101101110110000;
    rom_data[943]=16'b1000000101001100;
    rom_data[944]=16'b0101101111000111;
    rom_data[945]=16'b1000000001001101;
    rom_data[946]=16'b0101101111011110;
    rom_data[947]=16'b0111111101001000;
    rom_data[948]=16'b0101101111110101;
    rom_data[949]=16'b0111111000111101;
    rom_data[950]=16'b0101110000001100;
    rom_data[951]=16'b0111110100101101;
    rom_data[952]=16'b0101110000100010;
    rom_data[953]=16'b0111110000011000;
    rom_data[954]=16'b0101110000111000;
    rom_data[955]=16'b0111101011111111;
    rom_data[956]=16'b0101110001001110;
    rom_data[957]=16'b0111100111100001;
    rom_data[958]=16'b0101110001100100;
    rom_data[959]=16'b0111100011000000;
    rom_data[960]=16'b0101110001111010;
    rom_data[961]=16'b0111011110011011;
    rom_data[962]=16'b0101110010010000;
    rom_data[963]=16'b0111011001110010;
    rom_data[964]=16'b0101110010100101;
    rom_data[965]=16'b0111010101000111;
    rom_data[966]=16'b0101110010111011;
    rom_data[967]=16'b0111010000011000;
    rom_data[968]=16'b0101110011010000;
    rom_data[969]=16'b0111001011100111;
    rom_data[970]=16'b0101110011100101;
    rom_data[971]=16'b0111000110110100;
    rom_data[972]=16'b0101110011111010;
    rom_data[973]=16'b0111000001111110;
    rom_data[974]=16'b0101110100001111;
    rom_data[975]=16'b0110111101000111;
    rom_data[976]=16'b0101110100100100;
    rom_data[977]=16'b0110111000001101;
    rom_data[978]=16'b0101110100111001;
    rom_data[979]=16'b0110110011010010;
    rom_data[980]=16'b0101110101001110;
    rom_data[981]=16'b0110101110010110;
    rom_data[982]=16'b0101110101100011;
    rom_data[983]=16'b0110101001011000;
    rom_data[984]=16'b0101110101111000;
    rom_data[985]=16'b0110100100011000;
    rom_data[986]=16'b0101110110001100;
    rom_data[987]=16'b0110011111011000;
    rom_data[988]=16'b0101110110100001;
    rom_data[989]=16'b0110011010010111;
    rom_data[990]=16'b0101110110110110;
    rom_data[991]=16'b0110010101010101;
    rom_data[992]=16'b0101110111001010;
    rom_data[993]=16'b0110010000010010;
    rom_data[994]=16'b0101110111011111;
    rom_data[995]=16'b0110001011001111;
    rom_data[996]=16'b0101110111110100;
    rom_data[997]=16'b0110000110001011;
    rom_data[998]=16'b0101111000001000;
    rom_data[999]=16'b0110000001000111;
    rom_data[1000]=16'b0101111000011101;
    rom_data[1001]=16'b0101111100000011;
    rom_data[1002]=16'b0101111000110010;
    rom_data[1003]=16'b0101110110111111;
    rom_data[1004]=16'b0101111001000110;
    rom_data[1005]=16'b0101110001111011;
    rom_data[1006]=16'b0101111001011011;
    rom_data[1007]=16'b0101101100110111;
    rom_data[1008]=16'b0101111001110000;
    rom_data[1009]=16'b0101100111110011;
    rom_data[1010]=16'b0101111010000101;
    rom_data[1011]=16'b0101100010110000;
    rom_data[1012]=16'b0101111010011010;
    rom_data[1013]=16'b0101011101101101;
    rom_data[1014]=16'b0101111010101111;
    rom_data[1015]=16'b0101011000101011;
    rom_data[1016]=16'b0101111011000100;
    rom_data[1017]=16'b0101010011101010;
    rom_data[1018]=16'b0101111011011001;
    rom_data[1019]=16'b0101001110101010;
    rom_data[1020]=16'b0101111011101111;
    rom_data[1021]=16'b0101001001101011;
    rom_data[1022]=16'b0101111100000100;
    rom_data[1023]=16'b0101000100101100;
    rom_data[1024]=16'b0101111100011010;
    rom_data[1025]=16'b0100111111110000;
    rom_data[1026]=16'b0101111100101111;
    rom_data[1027]=16'b0100111010110100;
    rom_data[1028]=16'b0101111101000101;
    rom_data[1029]=16'b0100110101111011;
    rom_data[1030]=16'b0101111101011011;
    rom_data[1031]=16'b0100110001000011;
    rom_data[1032]=16'b0101111101110001;
    rom_data[1033]=16'b0100101100001101;
    rom_data[1034]=16'b0101111110000111;
    rom_data[1035]=16'b0100100111011001;
    rom_data[1036]=16'b0101111110011110;
    rom_data[1037]=16'b0100100010100111;
    rom_data[1038]=16'b0101111110110100;
    rom_data[1039]=16'b0100011101111000;
    rom_data[1040]=16'b0101111111001011;
    rom_data[1041]=16'b0100011001001100;
    rom_data[1042]=16'b0101111111100010;
    rom_data[1043]=16'b0100010100100010;
    rom_data[1044]=16'b0101111111111001;
    rom_data[1045]=16'b0100001111111100;
    rom_data[1046]=16'b0110000000010001;
    rom_data[1047]=16'b0100001011011001;
    rom_data[1048]=16'b0110000000101000;
    rom_data[1049]=16'b0100000110111001;
    rom_data[1050]=16'b0110000001000000;
    rom_data[1051]=16'b0100000010011110;
    rom_data[1052]=16'b0110000001011000;
    rom_data[1053]=16'b0011111110000111;
    rom_data[1054]=16'b0110000001110001;
    rom_data[1055]=16'b0011111001110100;
    rom_data[1056]=16'b0110000010001010;
    rom_data[1057]=16'b0011110101100110;
    rom_data[1058]=16'b0110000010100011;
    rom_data[1059]=16'b0011110001011101;
    rom_data[1060]=16'b0110000010111100;
    rom_data[1061]=16'b0011101101011010;
    rom_data[1062]=16'b0110000011010101;
    rom_data[1063]=16'b0011101001011101;
    rom_data[1064]=16'b0110000011101111;
    rom_data[1065]=16'b0011100101100110;
    rom_data[1066]=16'b0110000100001001;
    rom_data[1067]=16'b0011100001110110;
    rom_data[1068]=16'b0110000100100100;
    rom_data[1069]=16'b0011011110001110;
    rom_data[1070]=16'b0110000100111111;
    rom_data[1071]=16'b0011011010101101;
    rom_data[1072]=16'b0110000101011010;
    rom_data[1073]=16'b0011010111010101;
    rom_data[1074]=16'b0110000101110101;
    rom_data[1075]=16'b0011010100000110;
    rom_data[1076]=16'b0110000110010001;
    rom_data[1077]=16'b0011010001000001;
    rom_data[1078]=16'b0110000110101101;
    rom_data[1079]=16'b0011001110000110;
    rom_data[1080]=16'b0110000111001001;
    rom_data[1081]=16'b0011001011010110;
    rom_data[1082]=16'b0110000111100110;
    rom_data[1083]=16'b0011001000110010;
    rom_data[1084]=16'b0110001000000010;
    rom_data[1085]=16'b0011000110011010;
    rom_data[1086]=16'b0110001000011111;
    rom_data[1087]=16'b0011000100010000;
    rom_data[1088]=16'b0110001000111100;
    rom_data[1089]=16'b0011000010010011;
    rom_data[1090]=16'b0110001001011001;
    rom_data[1091]=16'b0011000000100101;
    rom_data[1092]=16'b0110001001110110;
    rom_data[1093]=16'b0010111111000110;
    rom_data[1094]=16'b0110001010010100;
    rom_data[1095]=16'b0010111101110110;
    rom_data[1096]=16'b0110001010110001;
    rom_data[1097]=16'b0010111100110111;
    rom_data[1098]=16'b0110001011001110;
    rom_data[1099]=16'b0010111100001001;
    rom_data[1100]=16'b0110001011101011;
    rom_data[1101]=16'b0010111011101100;
    rom_data[1102]=16'b0110001100001000;
    rom_data[1103]=16'b0010111011100000;
    rom_data[1104]=16'b0110001100100101;
    rom_data[1105]=16'b0010111011100110;
    rom_data[1106]=16'b0110001101000001;
    rom_data[1107]=16'b0010111011111101;
    rom_data[1108]=16'b0110001101011101;
    rom_data[1109]=16'b0010111100100110;
    rom_data[1110]=16'b0110001101111001;
    rom_data[1111]=16'b0010111101100000;
    rom_data[1112]=16'b0110001110010101;
    rom_data[1113]=16'b0010111110101010;
    rom_data[1114]=16'b0110001110110001;
    rom_data[1115]=16'b0011000000000101;
    rom_data[1116]=16'b0110001111001100;
    rom_data[1117]=16'b0011000001101111;
    rom_data[1118]=16'b0110001111100111;
    rom_data[1119]=16'b0011000011101001;
    rom_data[1120]=16'b0110010000000001;
    rom_data[1121]=16'b0011000101110001;
    rom_data[1122]=16'b0110010000011100;
    rom_data[1123]=16'b0011001000000110;
    rom_data[1124]=16'b0110010000110101;
    rom_data[1125]=16'b0011001010101001;
    rom_data[1126]=16'b0110010001001111;
    rom_data[1127]=16'b0011001101011000;
    rom_data[1128]=16'b0110010001101000;
    rom_data[1129]=16'b0011010000010010;
    rom_data[1130]=16'b0110010010000001;
    rom_data[1131]=16'b0011010011010111;
    rom_data[1132]=16'b0110010010011010;
    rom_data[1133]=16'b0011010110100111;
    rom_data[1134]=16'b0110010010110011;
    rom_data[1135]=16'b0011011001111111;
    rom_data[1136]=16'b0110010011001011;
    rom_data[1137]=16'b0011011101100001;
    rom_data[1138]=16'b0110010011100011;
    rom_data[1139]=16'b0011100001001010;
    rom_data[1140]=16'b0110010011111011;
    rom_data[1141]=16'b0011100100111100;
    rom_data[1142]=16'b0110010100010010;
    rom_data[1143]=16'b0011101000110100;
    rom_data[1144]=16'b0110010100101001;
    rom_data[1145]=16'b0011101100110011;
    rom_data[1146]=16'b0110010101000000;
    rom_data[1147]=16'b0011110000111000;
    rom_data[1148]=16'b0110010101010111;
    rom_data[1149]=16'b0011110101000011;
    rom_data[1150]=16'b0110010101101110;
    rom_data[1151]=16'b0011111001010011;
    rom_data[1152]=16'b0110010110000100;
    rom_data[1153]=16'b0011111101101000;
    rom_data[1154]=16'b0110010110011010;
    rom_data[1155]=16'b0100000010000001;
    rom_data[1156]=16'b0110010110110000;
    rom_data[1157]=16'b0100000110011111;
    rom_data[1158]=16'b0110010111000110;
    rom_data[1159]=16'b0100001011000000;
    rom_data[1160]=16'b0110010111011100;
    rom_data[1161]=16'b0100001111100101;
    rom_data[1162]=16'b0110010111110010;
    rom_data[1163]=16'b0100010100001110;
    rom_data[1164]=16'b0110011000000111;
    rom_data[1165]=16'b0100011000111001;
    rom_data[1166]=16'b0110011000011101;
    rom_data[1167]=16'b0100011101101000;
    rom_data[1168]=16'b0110011000110010;
    rom_data[1169]=16'b0100100010011001;
    rom_data[1170]=16'b0110011001000111;
    rom_data[1171]=16'b0100100111001100;
    rom_data[1172]=16'b0110011001011100;
    rom_data[1173]=16'b0100101100000010;
    rom_data[1174]=16'b0110011001110001;
    rom_data[1175]=16'b0100110000111001;
    rom_data[1176]=16'b0110011010000110;
    rom_data[1177]=16'b0100110101110011;
    rom_data[1178]=16'b0110011010011011;
    rom_data[1179]=16'b0100111010101110;
    rom_data[1180]=16'b0110011010110000;
    rom_data[1181]=16'b0100111111101011;
    rom_data[1182]=16'b0110011011000101;
    rom_data[1183]=16'b0101000100101001;
    rom_data[1184]=16'b0110011011011010;
    rom_data[1185]=16'b0101001001101000;
    rom_data[1186]=16'b0110011011101110;
    rom_data[1187]=16'b0101001110101000;
    rom_data[1188]=16'b0110011100000011;
    rom_data[1189]=16'b0101010011101001;
    rom_data[1190]=16'b0110011100011000;
    rom_data[1191]=16'b0101011000101011;
    rom_data[1192]=16'b0110011100101100;
    rom_data[1193]=16'b0101011101101110;
    rom_data[1194]=16'b0110011101000001;
    rom_data[1195]=16'b0101100010110001;
    rom_data[1196]=16'b0110011101010110;
    rom_data[1197]=16'b0101100111110101;
    rom_data[1198]=16'b0110011101101010;
    rom_data[1199]=16'b0101101100111001;
    rom_data[1200]=16'b0110011101111111;
    rom_data[1201]=16'b0101110001111101;
    rom_data[1202]=16'b0110011110010100;
    rom_data[1203]=16'b0101110111000001;
    rom_data[1204]=16'b0110011110101001;
    rom_data[1205]=16'b0101111100000101;
    rom_data[1206]=16'b0110011110111101;
    rom_data[1207]=16'b0110000001001001;
    rom_data[1208]=16'b0110011111010010;
    rom_data[1209]=16'b0110000110001101;
    rom_data[1210]=16'b0110011111100111;
    rom_data[1211]=16'b0110001011010000;
    rom_data[1212]=16'b0110011111111100;
    rom_data[1213]=16'b0110010000010011;
    rom_data[1214]=16'b0110100000010001;
    rom_data[1215]=16'b0110010101010101;
    rom_data[1216]=16'b0110100000100110;
    rom_data[1217]=16'b0110011010010110;
    rom_data[1218]=16'b0110100000111011;
    rom_data[1219]=16'b0110011111010110;
    rom_data[1220]=16'b0110100001010001;
    rom_data[1221]=16'b0110100100010110;
    rom_data[1222]=16'b0110100001100110;
    rom_data[1223]=16'b0110101001010100;
    rom_data[1224]=16'b0110100001111100;
    rom_data[1225]=16'b0110101110010000;
    rom_data[1226]=16'b0110100010010001;
    rom_data[1227]=16'b0110110011001100;
    rom_data[1228]=16'b0110100010100111;
    rom_data[1229]=16'b0110111000000110;
    rom_data[1230]=16'b0110100010111101;
    rom_data[1231]=16'b0110111100111101;
    rom_data[1232]=16'b0110100011010011;
    rom_data[1233]=16'b0111000001110011;
    rom_data[1234]=16'b0110100011101001;
    rom_data[1235]=16'b0111000110100111;
    rom_data[1236]=16'b0110100100000000;
    rom_data[1237]=16'b0111001011011001;
    rom_data[1238]=16'b0110100100010110;
    rom_data[1239]=16'b0111010000001000;
    rom_data[1240]=16'b0110100100101101;
    rom_data[1241]=16'b0111010100110100;
    rom_data[1242]=16'b0110100101000100;
    rom_data[1243]=16'b0111011001011110;
    rom_data[1244]=16'b0110100101011011;
    rom_data[1245]=16'b0111011110000100;
    rom_data[1246]=16'b0110100101110011;
    rom_data[1247]=16'b0111100010100111;
    rom_data[1248]=16'b0110100110001010;
    rom_data[1249]=16'b0111100111000111;
    rom_data[1250]=16'b0110100110100010;
    rom_data[1251]=16'b0111101011100010;
    rom_data[1252]=16'b0110100110111010;
    rom_data[1253]=16'b0111101111111010;
    rom_data[1254]=16'b0110100111010011;
    rom_data[1255]=16'b0111110100001100;
    rom_data[1256]=16'b0110100111101100;
    rom_data[1257]=16'b0111111000011010;
    rom_data[1258]=16'b0110101000000101;
    rom_data[1259]=16'b0111111100100011;
    rom_data[1260]=16'b0110101000011110;
    rom_data[1261]=16'b1000000000100110;
    rom_data[1262]=16'b0110101000110111;
    rom_data[1263]=16'b1000000100100011;
    rom_data[1264]=16'b0110101001010001;
    rom_data[1265]=16'b1000001000011010;
    rom_data[1266]=16'b0110101001101011;
    rom_data[1267]=16'b1000001100001010;
    rom_data[1268]=16'b0110101010000110;
    rom_data[1269]=16'b1000001111110010;
    rom_data[1270]=16'b0110101010100001;
    rom_data[1271]=16'b1000010011010011;
    rom_data[1272]=16'b0110101010111100;
    rom_data[1273]=16'b1000010110101011;
    rom_data[1274]=16'b0110101011010111;
    rom_data[1275]=16'b1000011001111010;
    rom_data[1276]=16'b0110101011110011;
    rom_data[1277]=16'b1000011100111111;
    rom_data[1278]=16'b0110101100001111;
    rom_data[1279]=16'b1000011111111010;
    rom_data[1280]=16'b0110101100101011;
    rom_data[1281]=16'b1000100010101010;
    rom_data[1282]=16'b0110101101001000;
    rom_data[1283]=16'b1000100101001110;
    rom_data[1284]=16'b0110101101100100;
    rom_data[1285]=16'b1000100111100110;
    rom_data[1286]=16'b0110101110000001;
    rom_data[1287]=16'b1000101001110000;
    rom_data[1288]=16'b0110101110011110;
    rom_data[1289]=16'b1000101011101101;
    rom_data[1290]=16'b0110101110111011;
    rom_data[1291]=16'b1000101101011011;
    rom_data[1292]=16'b0110101111011000;
    rom_data[1293]=16'b1000101110111011;
    rom_data[1294]=16'b0110101111110110;
    rom_data[1295]=16'b1000110000001010;
    rom_data[1296]=16'b0110110000010011;
    rom_data[1297]=16'b1000110001001001;
    rom_data[1298]=16'b0110110000110000;
    rom_data[1299]=16'b1000110001110111;
    rom_data[1300]=16'b0110110001001101;
    rom_data[1301]=16'b1000110010010100;
    rom_data[1302]=16'b0110110001101010;
    rom_data[1303]=16'b1000110010100000;
    rom_data[1304]=16'b0110110010000111;
    rom_data[1305]=16'b1000110010011010;
    rom_data[1306]=16'b0110110010100011;
    rom_data[1307]=16'b1000110010000011;
    rom_data[1308]=16'b0110110010111111;
    rom_data[1309]=16'b1000110001011010;
    rom_data[1310]=16'b0110110011011011;
    rom_data[1311]=16'b1000110000100000;
    rom_data[1312]=16'b0110110011110111;
    rom_data[1313]=16'b1000101111010110;
    rom_data[1314]=16'b0110110100010011;
    rom_data[1315]=16'b1000101101111011;
    rom_data[1316]=16'b0110110100101110;
    rom_data[1317]=16'b1000101100010001;
    rom_data[1318]=16'b0110110101001001;
    rom_data[1319]=16'b1000101010010111;
    rom_data[1320]=16'b0110110101100011;
    rom_data[1321]=16'b1000101000001111;
    rom_data[1322]=16'b0110110101111110;
    rom_data[1323]=16'b1000100101111010;
    rom_data[1324]=16'b0110110110011000;
    rom_data[1325]=16'b1000100011010111;
    rom_data[1326]=16'b0110110110110001;
    rom_data[1327]=16'b1000100000101000;
    rom_data[1328]=16'b0110110111001010;
    rom_data[1329]=16'b1000011101101110;
    rom_data[1330]=16'b0110110111100100;
    rom_data[1331]=16'b1000011010101001;
    rom_data[1332]=16'b0110110111111100;
    rom_data[1333]=16'b1000010111011001;
    rom_data[1334]=16'b0110111000010101;
    rom_data[1335]=16'b1000010100000001;
    rom_data[1336]=16'b0110111000101101;
    rom_data[1337]=16'b1000010000011111;
    rom_data[1338]=16'b0110111001000101;
    rom_data[1339]=16'b1000001100110101;
    rom_data[1340]=16'b0110111001011101;
    rom_data[1341]=16'b1000001001000100;
    rom_data[1342]=16'b0110111001110100;
    rom_data[1343]=16'b1000000101001100;
    rom_data[1344]=16'b0110111010001011;
    rom_data[1345]=16'b1000000001001101;
    rom_data[1346]=16'b0110111010100010;
    rom_data[1347]=16'b0111111101001000;
    rom_data[1348]=16'b0110111010111001;
    rom_data[1349]=16'b0111111000111101;
    rom_data[1350]=16'b0110111011010000;
    rom_data[1351]=16'b0111110100101101;
    rom_data[1352]=16'b0110111011100110;
    rom_data[1353]=16'b0111110000011000;
    rom_data[1354]=16'b0110111011111100;
    rom_data[1355]=16'b0111101011111111;
    rom_data[1356]=16'b0110111100010010;
    rom_data[1357]=16'b0111100111100001;
    rom_data[1358]=16'b0110111100101000;
    rom_data[1359]=16'b0111100010111111;
    rom_data[1360]=16'b0110111100111110;
    rom_data[1361]=16'b0111011110011010;
    rom_data[1362]=16'b0110111101010100;
    rom_data[1363]=16'b0111011001110010;
    rom_data[1364]=16'b0110111101101001;
    rom_data[1365]=16'b0111010101000110;
    rom_data[1366]=16'b0110111101111111;
    rom_data[1367]=16'b0111010000011000;
    rom_data[1368]=16'b0110111110010100;
    rom_data[1369]=16'b0111001011100111;
    rom_data[1370]=16'b0110111110101001;
    rom_data[1371]=16'b0111000110110100;
    rom_data[1372]=16'b0110111110111110;
    rom_data[1373]=16'b0111000001111110;
    rom_data[1374]=16'b0110111111010011;
    rom_data[1375]=16'b0110111101000110;
    rom_data[1376]=16'b0110111111101000;
    rom_data[1377]=16'b0110111000001101;
    rom_data[1378]=16'b0110111111111101;
    rom_data[1379]=16'b0110110011010010;
    rom_data[1380]=16'b0111000000010010;
    rom_data[1381]=16'b0110101110010101;
    rom_data[1382]=16'b0111000000100111;
    rom_data[1383]=16'b0110101001010111;
    rom_data[1384]=16'b0111000000111100;
    rom_data[1385]=16'b0110100100011000;
    rom_data[1386]=16'b0111000001010000;
    rom_data[1387]=16'b0110011111011000;
    rom_data[1388]=16'b0111000001100101;
    rom_data[1389]=16'b0110011010010110;
    rom_data[1390]=16'b0111000001111010;
    rom_data[1391]=16'b0110010101010100;
    rom_data[1392]=16'b0111000010001110;
    rom_data[1393]=16'b0110010000010010;
    rom_data[1394]=16'b0111000010100011;
    rom_data[1395]=16'b0110001011001111;
    rom_data[1396]=16'b0111000010111000;
    rom_data[1397]=16'b0110000110001011;
    rom_data[1398]=16'b0111000011001100;
    rom_data[1399]=16'b0110000001000111;
    rom_data[1400]=16'b0111000011100001;
    rom_data[1401]=16'b0101111100000011;
    rom_data[1402]=16'b0111000011110110;
    rom_data[1403]=16'b0101110110111111;
    rom_data[1404]=16'b0111000100001011;
    rom_data[1405]=16'b0101110001111011;
    rom_data[1406]=16'b0111000100011111;
    rom_data[1407]=16'b0101101100110111;
    rom_data[1408]=16'b0111000100110100;
    rom_data[1409]=16'b0101100111110011;
    rom_data[1410]=16'b0111000101001001;
    rom_data[1411]=16'b0101100010110000;
    rom_data[1412]=16'b0111000101011110;
    rom_data[1413]=16'b0101011101101101;
    rom_data[1414]=16'b0111000101110011;
    rom_data[1415]=16'b0101011000101011;
    rom_data[1416]=16'b0111000110001000;
    rom_data[1417]=16'b0101010011101010;
    rom_data[1418]=16'b0111000110011101;
    rom_data[1419]=16'b0101001110101001;
    rom_data[1420]=16'b0111000110110011;
    rom_data[1421]=16'b0101001001101010;
    rom_data[1422]=16'b0111000111001000;
    rom_data[1423]=16'b0101000100101100;
    rom_data[1424]=16'b0111000111011110;
    rom_data[1425]=16'b0100111111101111;
    rom_data[1426]=16'b0111000111110011;
    rom_data[1427]=16'b0100111010110100;
    rom_data[1428]=16'b0111001000001001;
    rom_data[1429]=16'b0100110101111010;
    rom_data[1430]=16'b0111001000011111;
    rom_data[1431]=16'b0100110001000010;
    rom_data[1432]=16'b0111001000110101;
    rom_data[1433]=16'b0100101100001100;
    rom_data[1434]=16'b0111001001001011;
    rom_data[1435]=16'b0100100111011000;
    rom_data[1436]=16'b0111001001100010;
    rom_data[1437]=16'b0100100010100111;
    rom_data[1438]=16'b0111001001111000;
    rom_data[1439]=16'b0100011101111000;
    rom_data[1440]=16'b0111001010001111;
    rom_data[1441]=16'b0100011001001011;
    rom_data[1442]=16'b0111001010100110;
    rom_data[1443]=16'b0100010100100010;
    rom_data[1444]=16'b0111001010111101;
    rom_data[1445]=16'b0100001111111011;
    rom_data[1446]=16'b0111001011010101;
    rom_data[1447]=16'b0100001011011000;
    rom_data[1448]=16'b0111001011101100;
    rom_data[1449]=16'b0100000110111001;
    rom_data[1450]=16'b0111001100000100;
    rom_data[1451]=16'b0100000010011110;
    rom_data[1452]=16'b0111001100011101;
    rom_data[1453]=16'b0011111110000110;
    rom_data[1454]=16'b0111001100110101;
    rom_data[1455]=16'b0011111001110011;
    rom_data[1456]=16'b0111001101001110;
    rom_data[1457]=16'b0011110101100110;
    rom_data[1458]=16'b0111001101100111;
    rom_data[1459]=16'b0011110001011101;
    rom_data[1460]=16'b0111001110000000;
    rom_data[1461]=16'b0011101101011010;
    rom_data[1462]=16'b0111001110011010;
    rom_data[1463]=16'b0011101001011101;
    rom_data[1464]=16'b0111001110110011;
    rom_data[1465]=16'b0011100101100110;
    rom_data[1466]=16'b0111001111001110;
    rom_data[1467]=16'b0011100001110110;
    rom_data[1468]=16'b0111001111101000;
    rom_data[1469]=16'b0011011110001110;
    rom_data[1470]=16'b0111010000000011;
    rom_data[1471]=16'b0011011010101101;
    rom_data[1472]=16'b0111010000011110;
    rom_data[1473]=16'b0011010111010101;
    rom_data[1474]=16'b0111010000111001;
    rom_data[1475]=16'b0011010100000110;
    rom_data[1476]=16'b0111010001010101;
    rom_data[1477]=16'b0011010001000001;
    rom_data[1478]=16'b0111010001110001;
    rom_data[1479]=16'b0011001110000110;
    rom_data[1480]=16'b0111010010001101;
    rom_data[1481]=16'b0011001011010110;
    rom_data[1482]=16'b0111010010101010;
    rom_data[1483]=16'b0011001000110010;
    rom_data[1484]=16'b0111010011000110;
    rom_data[1485]=16'b0011000110011010;
    rom_data[1486]=16'b0111010011100011;
    rom_data[1487]=16'b0011000100001111;
    rom_data[1488]=16'b0111010100000000;
    rom_data[1489]=16'b0011000010010011;
    rom_data[1490]=16'b0111010100011101;
    rom_data[1491]=16'b0011000000100100;
    rom_data[1492]=16'b0111010100111010;
    rom_data[1493]=16'b0010111111000101;
    rom_data[1494]=16'b0111010101011000;
    rom_data[1495]=16'b0010111101110110;
    rom_data[1496]=16'b0111010101110101;
    rom_data[1497]=16'b0010111100110111;
    rom_data[1498]=16'b0111010110010010;
    rom_data[1499]=16'b0010111100001001;
    rom_data[1500]=16'b0111010110101111;
    rom_data[1501]=16'b0010111011101100;
    rom_data[1502]=16'b0111010111001100;
    rom_data[1503]=16'b0010111011100000;
    rom_data[1504]=16'b0111010111101001;
    rom_data[1505]=16'b0010111011100110;
    rom_data[1506]=16'b0111011000000101;
    rom_data[1507]=16'b0010111011111101;
    rom_data[1508]=16'b0111011000100010;
    rom_data[1509]=16'b0010111100100110;
    rom_data[1510]=16'b0111011000111110;
    rom_data[1511]=16'b0010111101100000;
    rom_data[1512]=16'b0111011001011001;
    rom_data[1513]=16'b0010111110101010;
    rom_data[1514]=16'b0111011001110101;
    rom_data[1515]=16'b0011000000000101;
    rom_data[1516]=16'b0111011010010000;
    rom_data[1517]=16'b0011000001101111;
    rom_data[1518]=16'b0111011010101011;
    rom_data[1519]=16'b0011000011101001;
    rom_data[1520]=16'b0111011011000101;
    rom_data[1521]=16'b0011000101110001;
    rom_data[1522]=16'b0111011011100000;
    rom_data[1523]=16'b0011001000000111;
    rom_data[1524]=16'b0111011011111010;
    rom_data[1525]=16'b0011001010101001;
    rom_data[1526]=16'b0111011100010011;
    rom_data[1527]=16'b0011001101011000;
    rom_data[1528]=16'b0111011100101101;
    rom_data[1529]=16'b0011010000010010;
    rom_data[1530]=16'b0111011101000110;
    rom_data[1531]=16'b0011010011011000;
    rom_data[1532]=16'b0111011101011110;
    rom_data[1533]=16'b0011010110100111;
    rom_data[1534]=16'b0111011101110111;
    rom_data[1535]=16'b0011011010000000;
    rom_data[1536]=16'b0111011110001111;
    rom_data[1537]=16'b0011011101100001;
    rom_data[1538]=16'b0111011110100111;
    rom_data[1539]=16'b0011100001001011;
    rom_data[1540]=16'b0111011110111111;
    rom_data[1541]=16'b0011100100111100;
    rom_data[1542]=16'b0111011111010110;
    rom_data[1543]=16'b0011101000110100;
    rom_data[1544]=16'b0111011111101101;
    rom_data[1545]=16'b0011101100110011;
    rom_data[1546]=16'b0111100000000100;
    rom_data[1547]=16'b0011110000111000;
    rom_data[1548]=16'b0111100000011011;
    rom_data[1549]=16'b0011110101000011;
    rom_data[1550]=16'b0111100000110010;
    rom_data[1551]=16'b0011111001010011;
    rom_data[1552]=16'b0111100001001000;
    rom_data[1553]=16'b0011111101101000;
    rom_data[1554]=16'b0111100001011110;
    rom_data[1555]=16'b0100000010000010;
    rom_data[1556]=16'b0111100001110101;
    rom_data[1557]=16'b0100000110011111;
    rom_data[1558]=16'b0111100010001010;
    rom_data[1559]=16'b0100001011000001;
    rom_data[1560]=16'b0111100010100000;
    rom_data[1561]=16'b0100001111100110;
    rom_data[1562]=16'b0111100010110110;
    rom_data[1563]=16'b0100010100001110;
    rom_data[1564]=16'b0111100011001011;
    rom_data[1565]=16'b0100011000111010;
    rom_data[1566]=16'b0111100011100001;
    rom_data[1567]=16'b0100011101101000;
    rom_data[1568]=16'b0111100011110110;
    rom_data[1569]=16'b0100100010011001;
    rom_data[1570]=16'b0111100100001011;
    rom_data[1571]=16'b0100100111001101;
    rom_data[1572]=16'b0111100100100001;
    rom_data[1573]=16'b0100101100000010;
    rom_data[1574]=16'b0111100100110110;
    rom_data[1575]=16'b0100110000111010;
    rom_data[1576]=16'b0111100101001011;
    rom_data[1577]=16'b0100110101110011;
    rom_data[1578]=16'b0111100101011111;
    rom_data[1579]=16'b0100111010101110;
    rom_data[1580]=16'b0111100101110100;
    rom_data[1581]=16'b0100111111101011;
    rom_data[1582]=16'b0111100110001001;
    rom_data[1583]=16'b0101000100101001;
    rom_data[1584]=16'b0111100110011110;
    rom_data[1585]=16'b0101001001101000;
    rom_data[1586]=16'b0111100110110011;
    rom_data[1587]=16'b0101001110101000;
    rom_data[1588]=16'b0111100111000111;
    rom_data[1589]=16'b0101010011101010;
    rom_data[1590]=16'b0111100111011100;
    rom_data[1591]=16'b0101011000101100;
    rom_data[1592]=16'b0111100111110001;
    rom_data[1593]=16'b0101011101101110;
    rom_data[1594]=16'b0111101000000101;
    rom_data[1595]=16'b0101100010110010;
    rom_data[1596]=16'b0111101000011010;
    rom_data[1597]=16'b0101100111110101;
    rom_data[1598]=16'b0111101000101111;
    rom_data[1599]=16'b0101101100111001;
    rom_data[1600]=16'b0111101001000011;
    rom_data[1601]=16'b0101110001111101;
    rom_data[1602]=16'b0111101001011000;
    rom_data[1603]=16'b0101110111000001;
    rom_data[1604]=16'b0111101001101101;
    rom_data[1605]=16'b0101111100000110;
    rom_data[1606]=16'b0111101010000001;
    rom_data[1607]=16'b0110000001001010;
    rom_data[1608]=16'b0111101010010110;
    rom_data[1609]=16'b0110000110001101;
    rom_data[1610]=16'b0111101010101011;
    rom_data[1611]=16'b0110001011010000;
    rom_data[1612]=16'b0111101011000000;
    rom_data[1613]=16'b0110010000010011;
    rom_data[1614]=16'b0111101011010101;
    rom_data[1615]=16'b0110010101010101;
    rom_data[1616]=16'b0111101011101010;
    rom_data[1617]=16'b0110011010010110;
    rom_data[1618]=16'b0111101100000000;
    rom_data[1619]=16'b0110011111010111;
    rom_data[1620]=16'b0111101100010101;
    rom_data[1621]=16'b0110100100010110;
    rom_data[1622]=16'b0111101100101010;
    rom_data[1623]=16'b0110101001010100;
    rom_data[1624]=16'b0111101101000000;
    rom_data[1625]=16'b0110101110010001;
    rom_data[1626]=16'b0111101101010101;
    rom_data[1627]=16'b0110110011001100;
    rom_data[1628]=16'b0111101101101011;
    rom_data[1629]=16'b0110111000000110;
    rom_data[1630]=16'b0111101110000001;
    rom_data[1631]=16'b0110111100111110;
    rom_data[1632]=16'b0111101110010111;
    rom_data[1633]=16'b0111000001110100;
    rom_data[1634]=16'b0111101110101101;
    rom_data[1635]=16'b0111000110101000;
    rom_data[1636]=16'b0111101111000100;
    rom_data[1637]=16'b0111001011011001;
    rom_data[1638]=16'b0111101111011010;
    rom_data[1639]=16'b0111010000001000;
    rom_data[1640]=16'b0111101111110001;
    rom_data[1641]=16'b0111010100110101;
    rom_data[1642]=16'b0111110000001000;
    rom_data[1643]=16'b0111011001011110;
    rom_data[1644]=16'b0111110000011111;
    rom_data[1645]=16'b0111011110000101;
    rom_data[1646]=16'b0111110000110111;
    rom_data[1647]=16'b0111100010101000;
    rom_data[1648]=16'b0111110001001111;
    rom_data[1649]=16'b0111100111000111;
    rom_data[1650]=16'b0111110001100110;
    rom_data[1651]=16'b0111101011100011;
    rom_data[1652]=16'b0111110001111111;
    rom_data[1653]=16'b0111101111111010;
    rom_data[1654]=16'b0111110010010111;
    rom_data[1655]=16'b0111110100001101;
    rom_data[1656]=16'b0111110010110000;
    rom_data[1657]=16'b0111111000011011;
    rom_data[1658]=16'b0111110011001001;
    rom_data[1659]=16'b0111111100100011;
    rom_data[1660]=16'b0111110011100010;
    rom_data[1661]=16'b1000000000100110;
    rom_data[1662]=16'b0111110011111100;
    rom_data[1663]=16'b1000000100100100;
    rom_data[1664]=16'b0111110100010101;
    rom_data[1665]=16'b1000001000011010;
    rom_data[1666]=16'b0111110100110000;
    rom_data[1667]=16'b1000001100001010;
    rom_data[1668]=16'b0111110101001010;
    rom_data[1669]=16'b1000001111110011;
    rom_data[1670]=16'b0111110101100101;
    rom_data[1671]=16'b1000010011010011;
    rom_data[1672]=16'b0111110110000000;
    rom_data[1673]=16'b1000010110101011;
    rom_data[1674]=16'b0111110110011011;
    rom_data[1675]=16'b1000011001111010;
    rom_data[1676]=16'b0111110110110111;
    rom_data[1677]=16'b1000011100111111;
    rom_data[1678]=16'b0111110111010011;
    rom_data[1679]=16'b1000011111111010;
    rom_data[1680]=16'b0111110111101111;
    rom_data[1681]=16'b1000100010101010;
    rom_data[1682]=16'b0111111000001100;
    rom_data[1683]=16'b1000100101001110;
    rom_data[1684]=16'b0111111000101000;
    rom_data[1685]=16'b1000100111100110;
    rom_data[1686]=16'b0111111001000101;
    rom_data[1687]=16'b1000101001110001;
    rom_data[1688]=16'b0111111001100010;
    rom_data[1689]=16'b1000101011101101;
    rom_data[1690]=16'b0111111001111111;
    rom_data[1691]=16'b1000101101011100;
    rom_data[1692]=16'b0111111010011101;
    rom_data[1693]=16'b1000101110111011;
    rom_data[1694]=16'b0111111010111010;
    rom_data[1695]=16'b1000110000001010;
    rom_data[1696]=16'b0111111011010111;
    rom_data[1697]=16'b1000110001001001;
    rom_data[1698]=16'b0111111011110100;
    rom_data[1699]=16'b1000110001110111;
    rom_data[1700]=16'b0111111100010001;
    rom_data[1701]=16'b1000110010010100;
    rom_data[1702]=16'b0111111100101110;
    rom_data[1703]=16'b1000110010100000;
    rom_data[1704]=16'b0111111101001011;
    rom_data[1705]=16'b1000110010011010;
    rom_data[1706]=16'b0111111101100111;
    rom_data[1707]=16'b1000110010000011;
    rom_data[1708]=16'b0111111110000100;
    rom_data[1709]=16'b1000110001011010;
    rom_data[1710]=16'b0111111110100000;
    rom_data[1711]=16'b1000110000100000;
    rom_data[1712]=16'b0111111110111011;
    rom_data[1713]=16'b1000101111010110;
    rom_data[1714]=16'b0111111111010111;
    rom_data[1715]=16'b1000101101111011;
    rom_data[1716]=16'b0111111111110010;
    rom_data[1717]=16'b1000101100010001;
    rom_data[1718]=16'b1000000000001101;
    rom_data[1719]=16'b1000101010010111;
    rom_data[1720]=16'b1000000000100111;
    rom_data[1721]=16'b1000101000001111;
    rom_data[1722]=16'b1000000001000010;
    rom_data[1723]=16'b1000100101111001;
    rom_data[1724]=16'b1000000001011100;
    rom_data[1725]=16'b1000100011010111;
    rom_data[1726]=16'b1000000001110101;
    rom_data[1727]=16'b1000100000101000;
    rom_data[1728]=16'b1000000010001111;
    rom_data[1729]=16'b1000011101101101;
    rom_data[1730]=16'b1000000010101000;
    rom_data[1731]=16'b1000011010101000;
    rom_data[1732]=16'b1000000011000000;
    rom_data[1733]=16'b1000010111011001;
    rom_data[1734]=16'b1000000011011001;
    rom_data[1735]=16'b1000010100000000;
    rom_data[1736]=16'b1000000011110001;
    rom_data[1737]=16'b1000010000011111;
    rom_data[1738]=16'b1000000100001001;
    rom_data[1739]=16'b1000001100110101;
    rom_data[1740]=16'b1000000100100001;
    rom_data[1741]=16'b1000001001000100;
    rom_data[1742]=16'b1000000100111000;
    rom_data[1743]=16'b1000000101001011;
    rom_data[1744]=16'b1000000101001111;
    rom_data[1745]=16'b1000000001001101;
    rom_data[1746]=16'b1000000101100110;
    rom_data[1747]=16'b0111111101000111;
    rom_data[1748]=16'b1000000101111101;
    rom_data[1749]=16'b0111111000111101;
    rom_data[1750]=16'b1000000110010100;
    rom_data[1751]=16'b0111110100101101;
    rom_data[1752]=16'b1000000110101010;
    rom_data[1753]=16'b0111110000011000;
    rom_data[1754]=16'b1000000111000001;
    rom_data[1755]=16'b0111101011111110;
    rom_data[1756]=16'b1000000111010111;
    rom_data[1757]=16'b0111100111100001;
    rom_data[1758]=16'b1000000111101101;
    rom_data[1759]=16'b0111100010111111;
    rom_data[1760]=16'b1000001000000010;
    rom_data[1761]=16'b0111011110011010;
    rom_data[1762]=16'b1000001000011000;
    rom_data[1763]=16'b0111011001110010;
    rom_data[1764]=16'b1000001000101110;
    rom_data[1765]=16'b0111010101000110;
    rom_data[1766]=16'b1000001001000011;
    rom_data[1767]=16'b0111010000011000;
    rom_data[1768]=16'b1000001001011000;
    rom_data[1769]=16'b0111001011100111;
    rom_data[1770]=16'b1000001001101101;
    rom_data[1771]=16'b0111000110110011;
    rom_data[1772]=16'b1000001010000011;
    rom_data[1773]=16'b0111000001111110;
    rom_data[1774]=16'b1000001010011000;
    rom_data[1775]=16'b0110111101000110;
    rom_data[1776]=16'b1000001010101101;
    rom_data[1777]=16'b0110111000001101;
    rom_data[1778]=16'b1000001011000001;
    rom_data[1779]=16'b0110110011010001;
    rom_data[1780]=16'b1000001011010110;
    rom_data[1781]=16'b0110101110010101;
    rom_data[1782]=16'b1000001011101011;
    rom_data[1783]=16'b0110101001010111;
    rom_data[1784]=16'b1000001100000000;
    rom_data[1785]=16'b0110100100011000;
    rom_data[1786]=16'b1000001100010101;
    rom_data[1787]=16'b0110011111010111;
    rom_data[1788]=16'b1000001100101001;
    rom_data[1789]=16'b0110011010010110;
    rom_data[1790]=16'b1000001100111110;
    rom_data[1791]=16'b0110010101010100;
    rom_data[1792]=16'b1000001101010011;
    rom_data[1793]=16'b0110010000010001;
    rom_data[1794]=16'b1000001101100111;
    rom_data[1795]=16'b0110001011001110;
    rom_data[1796]=16'b1000001101111100;
    rom_data[1797]=16'b0110000110001011;
    rom_data[1798]=16'b1000001110010001;
    rom_data[1799]=16'b0110000001000111;
    rom_data[1800]=16'b1000001110100101;
    rom_data[1801]=16'b0101111100000011;
    rom_data[1802]=16'b1000001110111010;
    rom_data[1803]=16'b0101110110111110;
    rom_data[1804]=16'b1000001111001111;
    rom_data[1805]=16'b0101110001111010;
    rom_data[1806]=16'b1000001111100100;
    rom_data[1807]=16'b0101101100110110;
    rom_data[1808]=16'b1000001111111000;
    rom_data[1809]=16'b0101100111110011;
    rom_data[1810]=16'b1000010000001101;
    rom_data[1811]=16'b0101100010101111;
    rom_data[1812]=16'b1000010000100010;
    rom_data[1813]=16'b0101011101101101;
    rom_data[1814]=16'b1000010000110111;
    rom_data[1815]=16'b0101011000101011;
    rom_data[1816]=16'b1000010001001100;
    rom_data[1817]=16'b0101010011101001;
    rom_data[1818]=16'b1000010001100010;
    rom_data[1819]=16'b0101001110101001;
    rom_data[1820]=16'b1000010001110111;
    rom_data[1821]=16'b0101001001101010;
    rom_data[1822]=16'b1000010010001100;
    rom_data[1823]=16'b0101000100101100;
    rom_data[1824]=16'b1000010010100010;
    rom_data[1825]=16'b0100111111101111;
    rom_data[1826]=16'b1000010010110111;
    rom_data[1827]=16'b0100111010110100;
    rom_data[1828]=16'b1000010011001101;
    rom_data[1829]=16'b0100110101111010;
    rom_data[1830]=16'b1000010011100011;
    rom_data[1831]=16'b0100110001000010;
    rom_data[1832]=16'b1000010011111001;
    rom_data[1833]=16'b0100101100001100;
    rom_data[1834]=16'b1000010100010000;
    rom_data[1835]=16'b0100100111011000;
    rom_data[1836]=16'b1000010100100110;
    rom_data[1837]=16'b0100100010100111;
    rom_data[1838]=16'b1000010100111101;
    rom_data[1839]=16'b0100011101110111;
    rom_data[1840]=16'b1000010101010011;
    rom_data[1841]=16'b0100011001001011;
    rom_data[1842]=16'b1000010101101010;
    rom_data[1843]=16'b0100010100100010;
    rom_data[1844]=16'b1000010110000010;
    rom_data[1845]=16'b0100001111111011;
    rom_data[1846]=16'b1000010110011001;
    rom_data[1847]=16'b0100001011011000;
    rom_data[1848]=16'b1000010110110001;
    rom_data[1849]=16'b0100000110111001;
    rom_data[1850]=16'b1000010111001001;
    rom_data[1851]=16'b0100000010011101;
    rom_data[1852]=16'b1000010111100001;
    rom_data[1853]=16'b0011111110000110;
    rom_data[1854]=16'b1000010111111001;
    rom_data[1855]=16'b0011111001110011;
    rom_data[1856]=16'b1000011000010010;
    rom_data[1857]=16'b0011110101100101;
    rom_data[1858]=16'b1000011000101011;
    rom_data[1859]=16'b0011110001011101;
    rom_data[1860]=16'b1000011001000100;
    rom_data[1861]=16'b0011101101011001;
    rom_data[1862]=16'b1000011001011110;
    rom_data[1863]=16'b0011101001011100;
    rom_data[1864]=16'b1000011001111000;
    rom_data[1865]=16'b0011100101100110;
    rom_data[1866]=16'b1000011010010010;
    rom_data[1867]=16'b0011100001110110;
    rom_data[1868]=16'b1000011010101100;
    rom_data[1869]=16'b0011011110001101;
    rom_data[1870]=16'b1000011011000111;
    rom_data[1871]=16'b0011011010101101;
    rom_data[1872]=16'b1000011011100010;
    rom_data[1873]=16'b0011010111010101;
    rom_data[1874]=16'b1000011011111101;
    rom_data[1875]=16'b0011010100000110;
    rom_data[1876]=16'b1000011100011001;
    rom_data[1877]=16'b0011010001000001;
    rom_data[1878]=16'b1000011100110101;
    rom_data[1879]=16'b0011001110000110;
    rom_data[1880]=16'b1000011101010001;
    rom_data[1881]=16'b0011001011010110;
    rom_data[1882]=16'b1000011101101110;
    rom_data[1883]=16'b0011001000110010;
    rom_data[1884]=16'b1000011110001010;
    rom_data[1885]=16'b0011000110011010;
    rom_data[1886]=16'b1000011110100111;
    rom_data[1887]=16'b0011000100001111;
    rom_data[1888]=16'b1000011111000100;
    rom_data[1889]=16'b0011000010010011;
    rom_data[1890]=16'b1000011111100001;
    rom_data[1891]=16'b0011000000100100;
    rom_data[1892]=16'b1000011111111111;
    rom_data[1893]=16'b0010111111000101;
    rom_data[1894]=16'b1000100000011100;
    rom_data[1895]=16'b0010111101110110;
    rom_data[1896]=16'b1000100000111001;
    rom_data[1897]=16'b0010111100110111;
    rom_data[1898]=16'b1000100001010110;
    rom_data[1899]=16'b0010111100001001;
    rom_data[1900]=16'b1000100001110011;
    rom_data[1901]=16'b0010111011101100;
    rom_data[1902]=16'b1000100010010000;
    rom_data[1903]=16'b0010111011100000;
    rom_data[1904]=16'b1000100010101101;
    rom_data[1905]=16'b0010111011100110;
    rom_data[1906]=16'b1000100011001001;
    rom_data[1907]=16'b0010111011111101;
    rom_data[1908]=16'b1000100011100110;
    rom_data[1909]=16'b0010111100100110;
    rom_data[1910]=16'b1000100100000010;
    rom_data[1911]=16'b0010111101100000;
    rom_data[1912]=16'b1000100100011101;
    rom_data[1913]=16'b0010111110101010;
    rom_data[1914]=16'b1000100100111001;
    rom_data[1915]=16'b0011000000000101;
    rom_data[1916]=16'b1000100101010100;
    rom_data[1917]=16'b0011000001110000;
    rom_data[1918]=16'b1000100101101111;
    rom_data[1919]=16'b0011000011101001;
    rom_data[1920]=16'b1000100110001010;
    rom_data[1921]=16'b0011000101110001;
    rom_data[1922]=16'b1000100110100100;
    rom_data[1923]=16'b0011001000000111;
    rom_data[1924]=16'b1000100110111110;
    rom_data[1925]=16'b0011001010101001;
    rom_data[1926]=16'b1000100111010111;
    rom_data[1927]=16'b0011001101011000;
    rom_data[1928]=16'b1000100111110001;
    rom_data[1929]=16'b0011010000010011;
    rom_data[1930]=16'b1000101000001010;
    rom_data[1931]=16'b0011010011011000;
    rom_data[1932]=16'b1000101000100010;
    rom_data[1933]=16'b0011010110100111;
    rom_data[1934]=16'b1000101000111011;
    rom_data[1935]=16'b0011011010000000;
    rom_data[1936]=16'b1000101001010011;
    rom_data[1937]=16'b0011011101100001;
    rom_data[1938]=16'b1000101001101011;
    rom_data[1939]=16'b0011100001001011;
    rom_data[1940]=16'b1000101010000011;
    rom_data[1941]=16'b0011100100111100;
    rom_data[1942]=16'b1000101010011010;
    rom_data[1943]=16'b0011101000110101;
    rom_data[1944]=16'b1000101010110001;
    rom_data[1945]=16'b0011101100110100;
    rom_data[1946]=16'b1000101011001000;
    rom_data[1947]=16'b0011110000111001;
    rom_data[1948]=16'b1000101011011111;
    rom_data[1949]=16'b0011110101000011;
    rom_data[1950]=16'b1000101011110110;
    rom_data[1951]=16'b0011111001010100;
    rom_data[1952]=16'b1000101100001100;
    rom_data[1953]=16'b0011111101101000;
    rom_data[1954]=16'b1000101100100011;
    rom_data[1955]=16'b0100000010000010;
    rom_data[1956]=16'b1000101100111001;
    rom_data[1957]=16'b0100000110100000;
    rom_data[1958]=16'b1000101101001111;
    rom_data[1959]=16'b0100001011000001;
    rom_data[1960]=16'b1000101101100100;
    rom_data[1961]=16'b0100001111100110;
    rom_data[1962]=16'b1000101101111010;
    rom_data[1963]=16'b0100010100001111;
    rom_data[1964]=16'b1000101110010000;
    rom_data[1965]=16'b0100011000111010;
    rom_data[1966]=16'b1000101110100101;
    rom_data[1967]=16'b0100011101101001;
    rom_data[1968]=16'b1000101110111010;
    rom_data[1969]=16'b0100100010011010;
    rom_data[1970]=16'b1000101111010000;
    rom_data[1971]=16'b0100100111001101;
    rom_data[1972]=16'b1000101111100101;
    rom_data[1973]=16'b0100101100000011;
    rom_data[1974]=16'b1000101111111010;
    rom_data[1975]=16'b0100110000111010;
    rom_data[1976]=16'b1000110000001111;
    rom_data[1977]=16'b0100110101110100;
    rom_data[1978]=16'b1000110000100100;
    rom_data[1979]=16'b0100111010101111;
    rom_data[1980]=16'b1000110000111000;
    rom_data[1981]=16'b0100111111101011;
    rom_data[1982]=16'b1000110001001101;
    rom_data[1983]=16'b0101000100101001;
    rom_data[1984]=16'b1000110001100010;
    rom_data[1985]=16'b0101001001101001;
    rom_data[1986]=16'b1000110001110111;
    rom_data[1987]=16'b0101001110101001;
    rom_data[1988]=16'b1000110010001011;
    rom_data[1989]=16'b0101010011101010;
    rom_data[1990]=16'b1000110010100000;
    rom_data[1991]=16'b0101011000101100;
    rom_data[1992]=16'b1000110010100000;
    rom_data[1993]=16'b0101011101101111;
    rom_data[1994]=16'b1000110010001011;
    rom_data[1995]=16'b0101100010110010;
    rom_data[1996]=16'b1000110001110111;
    rom_data[1997]=16'b0101100111110110;
    rom_data[1998]=16'b1000110001100010;
    rom_data[1999]=16'b0101101100111010;
    rom_data[2000]=16'b1000110001001101;
    rom_data[2001]=16'b0101110001111110;
    rom_data[2002]=16'b1000110000111000;
    rom_data[2003]=16'b0101110111000010;
    rom_data[2004]=16'b1000110000100100;
    rom_data[2005]=16'b0101111100000110;
    rom_data[2006]=16'b1000110000001111;
    rom_data[2007]=16'b0110000001001010;
    rom_data[2008]=16'b1000101111111010;
    rom_data[2009]=16'b0110000110001110;
    rom_data[2010]=16'b1000101111100101;
    rom_data[2011]=16'b0110001011010001;
    rom_data[2012]=16'b1000101111010000;
    rom_data[2013]=16'b0110010000010011;
    rom_data[2014]=16'b1000101110111010;
    rom_data[2015]=16'b0110010101010101;
    rom_data[2016]=16'b1000101110100101;
    rom_data[2017]=16'b0110011010010111;
    rom_data[2018]=16'b1000101110010000;
    rom_data[2019]=16'b0110011111010111;
    rom_data[2020]=16'b1000101101111010;
    rom_data[2021]=16'b0110100100010110;
    rom_data[2022]=16'b1000101101100100;
    rom_data[2023]=16'b0110101001010100;
    rom_data[2024]=16'b1000101101001111;
    rom_data[2025]=16'b0110101110010001;
    rom_data[2026]=16'b1000101100111001;
    rom_data[2027]=16'b0110110011001101;
    rom_data[2028]=16'b1000101100100011;
    rom_data[2029]=16'b0110111000000110;
    rom_data[2030]=16'b1000101100001100;
    rom_data[2031]=16'b0110111100111110;
    rom_data[2032]=16'b1000101011110110;
    rom_data[2033]=16'b0111000001110100;
    rom_data[2034]=16'b1000101011011111;
    rom_data[2035]=16'b0111000110101000;
    rom_data[2036]=16'b1000101011001000;
    rom_data[2037]=16'b0111001011011010;
    rom_data[2038]=16'b1000101010110001;
    rom_data[2039]=16'b0111010000001001;
    rom_data[2040]=16'b1000101010011010;
    rom_data[2041]=16'b0111010100110101;
    rom_data[2042]=16'b1000101010000011;
    rom_data[2043]=16'b0111011001011111;
    rom_data[2044]=16'b1000101001101011;
    rom_data[2045]=16'b0111011110000101;
    rom_data[2046]=16'b1000101001010011;
    rom_data[2047]=16'b0111100010101000;
    rom_data[2048]=16'b1000101000111011;
    rom_data[2049]=16'b0111100111000111;
    rom_data[2050]=16'b1000101000100010;
    rom_data[2051]=16'b0111101011100011;
    rom_data[2052]=16'b1000101000001010;
    rom_data[2053]=16'b0111101111111010;
    rom_data[2054]=16'b1000100111110001;
    rom_data[2055]=16'b0111110100001101;
    rom_data[2056]=16'b1000100111010111;
    rom_data[2057]=16'b0111111000011011;
    rom_data[2058]=16'b1000100110111110;
    rom_data[2059]=16'b0111111100100100;
    rom_data[2060]=16'b1000100110100100;
    rom_data[2061]=16'b1000000000100111;
    rom_data[2062]=16'b1000100110001010;
    rom_data[2063]=16'b1000000100100100;
    rom_data[2064]=16'b1000100101101111;
    rom_data[2065]=16'b1000001000011011;
    rom_data[2066]=16'b1000100101010100;
    rom_data[2067]=16'b1000001100001010;
    rom_data[2068]=16'b1000100100111001;
    rom_data[2069]=16'b1000001111110011;
    rom_data[2070]=16'b1000100100011101;
    rom_data[2071]=16'b1000010011010011;
    rom_data[2072]=16'b1000100100000010;
    rom_data[2073]=16'b1000010110101011;
    rom_data[2074]=16'b1000100011100110;
    rom_data[2075]=16'b1000011001111010;
    rom_data[2076]=16'b1000100011001001;
    rom_data[2077]=16'b1000011101000000;
    rom_data[2078]=16'b1000100010101101;
    rom_data[2079]=16'b1000011111111010;
    rom_data[2080]=16'b1000100010010000;
    rom_data[2081]=16'b1000100010101010;
    rom_data[2082]=16'b1000100001110011;
    rom_data[2083]=16'b1000100101001110;
    rom_data[2084]=16'b1000100001010110;
    rom_data[2085]=16'b1000100111100110;
    rom_data[2086]=16'b1000100000111001;
    rom_data[2087]=16'b1000101001110001;
    rom_data[2088]=16'b1000100000011100;
    rom_data[2089]=16'b1000101011101101;
    rom_data[2090]=16'b1000011111111111;
    rom_data[2091]=16'b1000101101011100;
    rom_data[2092]=16'b1000011111100001;
    rom_data[2093]=16'b1000101110111011;
    rom_data[2094]=16'b1000011111000100;
    rom_data[2095]=16'b1000110000001010;
    rom_data[2096]=16'b1000011110100111;
    rom_data[2097]=16'b1000110001001001;
    rom_data[2098]=16'b1000011110001010;
    rom_data[2099]=16'b1000110001110111;
    rom_data[2100]=16'b1000011101101110;
    rom_data[2101]=16'b1000110010010100;
    rom_data[2102]=16'b1000011101010001;
    rom_data[2103]=16'b1000110010100000;
    rom_data[2104]=16'b1000011100110101;
    rom_data[2105]=16'b1000110010011010;
    rom_data[2106]=16'b1000011100011001;
    rom_data[2107]=16'b1000110010000011;
    rom_data[2108]=16'b1000011011111101;
    rom_data[2109]=16'b1000110001011010;
    rom_data[2110]=16'b1000011011100010;
    rom_data[2111]=16'b1000110000100000;
    rom_data[2112]=16'b1000011011000111;
    rom_data[2113]=16'b1000101111010110;
    rom_data[2114]=16'b1000011010101100;
    rom_data[2115]=16'b1000101101111011;
    rom_data[2116]=16'b1000011010010010;
    rom_data[2117]=16'b1000101100010000;
    rom_data[2118]=16'b1000011001111000;
    rom_data[2119]=16'b1000101010010111;
    rom_data[2120]=16'b1000011001011110;
    rom_data[2121]=16'b1000101000001111;
    rom_data[2122]=16'b1000011001000100;
    rom_data[2123]=16'b1000100101111001;
    rom_data[2124]=16'b1000011000101011;
    rom_data[2125]=16'b1000100011010111;
    rom_data[2126]=16'b1000011000010010;
    rom_data[2127]=16'b1000100000101000;
    rom_data[2128]=16'b1000010111111001;
    rom_data[2129]=16'b1000011101101101;
    rom_data[2130]=16'b1000010111100001;
    rom_data[2131]=16'b1000011010101000;
    rom_data[2132]=16'b1000010111001001;
    rom_data[2133]=16'b1000010111011001;
    rom_data[2134]=16'b1000010110110001;
    rom_data[2135]=16'b1000010100000000;
    rom_data[2136]=16'b1000010110011001;
    rom_data[2137]=16'b1000010000011111;
    rom_data[2138]=16'b1000010110000010;
    rom_data[2139]=16'b1000001100110101;
    rom_data[2140]=16'b1000010101101010;
    rom_data[2141]=16'b1000001001000100;
    rom_data[2142]=16'b1000010101010011;
    rom_data[2143]=16'b1000000101001011;
    rom_data[2144]=16'b1000010100111101;
    rom_data[2145]=16'b1000000001001100;
    rom_data[2146]=16'b1000010100100110;
    rom_data[2147]=16'b0111111101000111;
    rom_data[2148]=16'b1000010100010000;
    rom_data[2149]=16'b0111111000111100;
    rom_data[2150]=16'b1000010011111001;
    rom_data[2151]=16'b0111110100101100;
    rom_data[2152]=16'b1000010011100011;
    rom_data[2153]=16'b0111110000010111;
    rom_data[2154]=16'b1000010011001101;
    rom_data[2155]=16'b0111101011111110;
    rom_data[2156]=16'b1000010010110111;
    rom_data[2157]=16'b0111100111100000;
    rom_data[2158]=16'b1000010010100010;
    rom_data[2159]=16'b0111100010111111;
    rom_data[2160]=16'b1000010010001100;
    rom_data[2161]=16'b0111011110011010;
    rom_data[2162]=16'b1000010001110111;
    rom_data[2163]=16'b0111011001110001;
    rom_data[2164]=16'b1000010001100010;
    rom_data[2165]=16'b0111010101000110;
    rom_data[2166]=16'b1000010001001100;
    rom_data[2167]=16'b0111010000010111;
    rom_data[2168]=16'b1000010000110111;
    rom_data[2169]=16'b0111001011100110;
    rom_data[2170]=16'b1000010000100010;
    rom_data[2171]=16'b0111000110110011;
    rom_data[2172]=16'b1000010000001101;
    rom_data[2173]=16'b0111000001111101;
    rom_data[2174]=16'b1000001111111000;
    rom_data[2175]=16'b0110111101000110;
    rom_data[2176]=16'b1000001111100100;
    rom_data[2177]=16'b0110111000001100;
    rom_data[2178]=16'b1000001111001111;
    rom_data[2179]=16'b0110110011010001;
    rom_data[2180]=16'b1000001110111010;
    rom_data[2181]=16'b0110101110010100;
    rom_data[2182]=16'b1000001110100101;
    rom_data[2183]=16'b0110101001010110;
    rom_data[2184]=16'b1000001110010001;
    rom_data[2185]=16'b0110100100010111;
    rom_data[2186]=16'b1000001101111100;
    rom_data[2187]=16'b0110011111010111;
    rom_data[2188]=16'b1000001101100111;
    rom_data[2189]=16'b0110011010010110;
    rom_data[2190]=16'b1000001101010011;
    rom_data[2191]=16'b0110010101010100;
    rom_data[2192]=16'b1000001100111110;
    rom_data[2193]=16'b0110010000010001;
    rom_data[2194]=16'b1000001100101001;
    rom_data[2195]=16'b0110001011001110;
    rom_data[2196]=16'b1000001100010101;
    rom_data[2197]=16'b0110000110001010;
    rom_data[2198]=16'b1000001100000000;
    rom_data[2199]=16'b0110000001000110;
    rom_data[2200]=16'b1000001011101011;
    rom_data[2201]=16'b0101111100000010;
    rom_data[2202]=16'b1000001011010110;
    rom_data[2203]=16'b0101110110111110;
    rom_data[2204]=16'b1000001011000001;
    rom_data[2205]=16'b0101110001111010;
    rom_data[2206]=16'b1000001010101101;
    rom_data[2207]=16'b0101101100110110;
    rom_data[2208]=16'b1000001010011000;
    rom_data[2209]=16'b0101100111110010;
    rom_data[2210]=16'b1000001010000011;
    rom_data[2211]=16'b0101100010101111;
    rom_data[2212]=16'b1000001001101101;
    rom_data[2213]=16'b0101011101101100;
    rom_data[2214]=16'b1000001001011000;
    rom_data[2215]=16'b0101011000101010;
    rom_data[2216]=16'b1000001001000011;
    rom_data[2217]=16'b0101010011101001;
    rom_data[2218]=16'b1000001000101110;
    rom_data[2219]=16'b0101001110101001;
    rom_data[2220]=16'b1000001000011000;
    rom_data[2221]=16'b0101001001101001;
    rom_data[2222]=16'b1000001000000010;
    rom_data[2223]=16'b0101000100101011;
    rom_data[2224]=16'b1000000111101101;
    rom_data[2225]=16'b0100111111101111;
    rom_data[2226]=16'b1000000111010111;
    rom_data[2227]=16'b0100111010110011;
    rom_data[2228]=16'b1000000111000001;
    rom_data[2229]=16'b0100110101111010;
    rom_data[2230]=16'b1000000110101010;
    rom_data[2231]=16'b0100110001000010;
    rom_data[2232]=16'b1000000110010100;
    rom_data[2233]=16'b0100101100001100;
    rom_data[2234]=16'b1000000101111101;
    rom_data[2235]=16'b0100100111011000;
    rom_data[2236]=16'b1000000101100110;
    rom_data[2237]=16'b0100100010100110;
    rom_data[2238]=16'b1000000101001111;
    rom_data[2239]=16'b0100011101110111;
    rom_data[2240]=16'b1000000100111000;
    rom_data[2241]=16'b0100011001001011;
    rom_data[2242]=16'b1000000100100001;
    rom_data[2243]=16'b0100010100100001;
    rom_data[2244]=16'b1000000100001001;
    rom_data[2245]=16'b0100001111111011;
    rom_data[2246]=16'b1000000011110001;
    rom_data[2247]=16'b0100001011011000;
    rom_data[2248]=16'b1000000011011001;
    rom_data[2249]=16'b0100000110111000;
    rom_data[2250]=16'b1000000011000000;
    rom_data[2251]=16'b0100000010011101;
    rom_data[2252]=16'b1000000010101000;
    rom_data[2253]=16'b0011111110000110;
    rom_data[2254]=16'b1000000010001111;
    rom_data[2255]=16'b0011111001110011;
    rom_data[2256]=16'b1000000001110101;
    rom_data[2257]=16'b0011110101100101;
    rom_data[2258]=16'b1000000001011100;
    rom_data[2259]=16'b0011110001011100;
    rom_data[2260]=16'b1000000001000010;
    rom_data[2261]=16'b0011101101011001;
    rom_data[2262]=16'b1000000000100111;
    rom_data[2263]=16'b0011101001011100;
    rom_data[2264]=16'b1000000000001101;
    rom_data[2265]=16'b0011100101100101;
    rom_data[2266]=16'b0111111111110010;
    rom_data[2267]=16'b0011100001110101;
    rom_data[2268]=16'b0111111111010111;
    rom_data[2269]=16'b0011011110001101;
    rom_data[2270]=16'b0111111110111011;
    rom_data[2271]=16'b0011011010101101;
    rom_data[2272]=16'b0111111110100000;
    rom_data[2273]=16'b0011010111010101;
    rom_data[2274]=16'b0111111110000100;
    rom_data[2275]=16'b0011010100000110;
    rom_data[2276]=16'b0111111101100111;
    rom_data[2277]=16'b0011010001000000;
    rom_data[2278]=16'b0111111101001011;
    rom_data[2279]=16'b0011001110000101;
    rom_data[2280]=16'b0111111100101110;
    rom_data[2281]=16'b0011001011010110;
    rom_data[2282]=16'b0111111100010001;
    rom_data[2283]=16'b0011001000110001;
    rom_data[2284]=16'b0111111011110100;
    rom_data[2285]=16'b0011000110011010;
    rom_data[2286]=16'b0111111011010111;
    rom_data[2287]=16'b0011000100001111;
    rom_data[2288]=16'b0111111010111010;
    rom_data[2289]=16'b0011000010010010;
    rom_data[2290]=16'b0111111010011101;
    rom_data[2291]=16'b0011000000100100;
    rom_data[2292]=16'b0111111001111111;
    rom_data[2293]=16'b0010111111000101;
    rom_data[2294]=16'b0111111001100010;
    rom_data[2295]=16'b0010111101110110;
    rom_data[2296]=16'b0111111001000101;
    rom_data[2297]=16'b0010111100110111;
    rom_data[2298]=16'b0111111000101000;
    rom_data[2299]=16'b0010111100001001;
    rom_data[2300]=16'b0111111000001100;
    rom_data[2301]=16'b0010111011101100;
    rom_data[2302]=16'b0111110111101111;
    rom_data[2303]=16'b0010111011100000;
    rom_data[2304]=16'b0111110111010011;
    rom_data[2305]=16'b0010111011100110;
    rom_data[2306]=16'b0111110110110111;
    rom_data[2307]=16'b0010111011111101;
    rom_data[2308]=16'b0111110110011011;
    rom_data[2309]=16'b0010111100100110;
    rom_data[2310]=16'b0111110110000000;
    rom_data[2311]=16'b0010111101100000;
    rom_data[2312]=16'b0111110101100101;
    rom_data[2313]=16'b0010111110101010;
    rom_data[2314]=16'b0111110101001010;
    rom_data[2315]=16'b0011000000000101;
    rom_data[2316]=16'b0111110100110000;
    rom_data[2317]=16'b0011000001110000;
    rom_data[2318]=16'b0111110100010101;
    rom_data[2319]=16'b0011000011101001;
    rom_data[2320]=16'b0111110011111100;
    rom_data[2321]=16'b0011000101110001;
    rom_data[2322]=16'b0111110011100010;
    rom_data[2323]=16'b0011001000000111;
    rom_data[2324]=16'b0111110011001001;
    rom_data[2325]=16'b0011001010101010;
    rom_data[2326]=16'b0111110010110000;
    rom_data[2327]=16'b0011001101011000;
    rom_data[2328]=16'b0111110010010111;
    rom_data[2329]=16'b0011010000010011;
    rom_data[2330]=16'b0111110001111111;
    rom_data[2331]=16'b0011010011011000;
    rom_data[2332]=16'b0111110001100110;
    rom_data[2333]=16'b0011010110100111;
    rom_data[2334]=16'b0111110001001111;
    rom_data[2335]=16'b0011011010000000;
    rom_data[2336]=16'b0111110000110111;
    rom_data[2337]=16'b0011011101100010;
    rom_data[2338]=16'b0111110000011111;
    rom_data[2339]=16'b0011100001001011;
    rom_data[2340]=16'b0111110000001000;
    rom_data[2341]=16'b0011100100111101;
    rom_data[2342]=16'b0111101111110001;
    rom_data[2343]=16'b0011101000110101;
    rom_data[2344]=16'b0111101111011010;
    rom_data[2345]=16'b0011101100110100;
    rom_data[2346]=16'b0111101111000100;
    rom_data[2347]=16'b0011110000111001;
    rom_data[2348]=16'b0111101110101101;
    rom_data[2349]=16'b0011110101000100;
    rom_data[2350]=16'b0111101110010111;
    rom_data[2351]=16'b0011111001010100;
    rom_data[2352]=16'b0111101110000001;
    rom_data[2353]=16'b0011111101101001;
    rom_data[2354]=16'b0111101101101011;
    rom_data[2355]=16'b0100000010000010;
    rom_data[2356]=16'b0111101101010101;
    rom_data[2357]=16'b0100000110100000;
    rom_data[2358]=16'b0111101101000000;
    rom_data[2359]=16'b0100001011000001;
    rom_data[2360]=16'b0111101100101010;
    rom_data[2361]=16'b0100001111100111;
    rom_data[2362]=16'b0111101100010101;
    rom_data[2363]=16'b0100010100001111;
    rom_data[2364]=16'b0111101100000000;
    rom_data[2365]=16'b0100011000111011;
    rom_data[2366]=16'b0111101011101010;
    rom_data[2367]=16'b0100011101101001;
    rom_data[2368]=16'b0111101011010101;
    rom_data[2369]=16'b0100100010011010;
    rom_data[2370]=16'b0111101011000000;
    rom_data[2371]=16'b0100100111001101;
    rom_data[2372]=16'b0111101010101011;
    rom_data[2373]=16'b0100101100000011;
    rom_data[2374]=16'b0111101010010110;
    rom_data[2375]=16'b0100110000111010;
    rom_data[2376]=16'b0111101010000001;
    rom_data[2377]=16'b0100110101110100;
    rom_data[2378]=16'b0111101001101101;
    rom_data[2379]=16'b0100111010101111;
    rom_data[2380]=16'b0111101001011000;
    rom_data[2381]=16'b0100111111101100;
    rom_data[2382]=16'b0111101001000011;
    rom_data[2383]=16'b0101000100101010;
    rom_data[2384]=16'b0111101000101111;
    rom_data[2385]=16'b0101001001101001;
    rom_data[2386]=16'b0111101000011010;
    rom_data[2387]=16'b0101001110101001;
    rom_data[2388]=16'b0111101000000101;
    rom_data[2389]=16'b0101010011101010;
    rom_data[2390]=16'b0111100111110001;
    rom_data[2391]=16'b0101011000101100;
    rom_data[2392]=16'b0111100111011100;
    rom_data[2393]=16'b0101011101101111;
    rom_data[2394]=16'b0111100111000111;
    rom_data[2395]=16'b0101100010110010;
    rom_data[2396]=16'b0111100110110011;
    rom_data[2397]=16'b0101100111110110;
    rom_data[2398]=16'b0111100110011110;
    rom_data[2399]=16'b0101101100111010;
    rom_data[2400]=16'b0111100110001001;
    rom_data[2401]=16'b0101110001111110;
    rom_data[2402]=16'b0111100101110100;
    rom_data[2403]=16'b0101110111000010;
    rom_data[2404]=16'b0111100101011111;
    rom_data[2405]=16'b0101111100000110;
    rom_data[2406]=16'b0111100101001011;
    rom_data[2407]=16'b0110000001001010;
    rom_data[2408]=16'b0111100100110110;
    rom_data[2409]=16'b0110000110001110;
    rom_data[2410]=16'b0111100100100001;
    rom_data[2411]=16'b0110001011010001;
    rom_data[2412]=16'b0111100100001011;
    rom_data[2413]=16'b0110010000010100;
    rom_data[2414]=16'b0111100011110110;
    rom_data[2415]=16'b0110010101010110;
    rom_data[2416]=16'b0111100011100001;
    rom_data[2417]=16'b0110011010010111;
    rom_data[2418]=16'b0111100011001011;
    rom_data[2419]=16'b0110011111010111;
    rom_data[2420]=16'b0111100010110110;
    rom_data[2421]=16'b0110100100010111;
    rom_data[2422]=16'b0111100010100000;
    rom_data[2423]=16'b0110101001010101;
    rom_data[2424]=16'b0111100010001010;
    rom_data[2425]=16'b0110101110010010;
    rom_data[2426]=16'b0111100001110101;
    rom_data[2427]=16'b0110110011001101;
    rom_data[2428]=16'b0111100001011110;
    rom_data[2429]=16'b0110111000000111;
    rom_data[2430]=16'b0111100001001000;
    rom_data[2431]=16'b0110111100111111;
    rom_data[2432]=16'b0111100000110010;
    rom_data[2433]=16'b0111000001110101;
    rom_data[2434]=16'b0111100000011011;
    rom_data[2435]=16'b0111000110101000;
    rom_data[2436]=16'b0111100000000100;
    rom_data[2437]=16'b0111001011011010;
    rom_data[2438]=16'b0111011111101101;
    rom_data[2439]=16'b0111010000001001;
    rom_data[2440]=16'b0111011111010110;
    rom_data[2441]=16'b0111010100110101;
    rom_data[2442]=16'b0111011110111111;
    rom_data[2443]=16'b0111011001011111;
    rom_data[2444]=16'b0111011110100111;
    rom_data[2445]=16'b0111011110000101;
    rom_data[2446]=16'b0111011110001111;
    rom_data[2447]=16'b0111100010101000;
    rom_data[2448]=16'b0111011101110111;
    rom_data[2449]=16'b0111100111001000;
    rom_data[2450]=16'b0111011101011110;
    rom_data[2451]=16'b0111101011100011;
    rom_data[2452]=16'b0111011101000110;
    rom_data[2453]=16'b0111101111111011;
    rom_data[2454]=16'b0111011100101101;
    rom_data[2455]=16'b0111110100001101;
    rom_data[2456]=16'b0111011100010011;
    rom_data[2457]=16'b0111111000011011;
    rom_data[2458]=16'b0111011011111010;
    rom_data[2459]=16'b0111111100100100;
    rom_data[2460]=16'b0111011011100000;
    rom_data[2461]=16'b1000000000100111;
    rom_data[2462]=16'b0111011011000101;
    rom_data[2463]=16'b1000000100100100;
    rom_data[2464]=16'b0111011010101011;
    rom_data[2465]=16'b1000001000011011;
    rom_data[2466]=16'b0111011010010000;
    rom_data[2467]=16'b1000001100001011;
    rom_data[2468]=16'b0111011001110101;
    rom_data[2469]=16'b1000001111110011;
    rom_data[2470]=16'b0111011001011001;
    rom_data[2471]=16'b1000010011010100;
    rom_data[2472]=16'b0111011000111110;
    rom_data[2473]=16'b1000010110101100;
    rom_data[2474]=16'b0111011000100010;
    rom_data[2475]=16'b1000011001111011;
    rom_data[2476]=16'b0111011000000101;
    rom_data[2477]=16'b1000011101000000;
    rom_data[2478]=16'b0111010111101001;
    rom_data[2479]=16'b1000011111111011;
    rom_data[2480]=16'b0111010111001100;
    rom_data[2481]=16'b1000100010101010;
    rom_data[2482]=16'b0111010110101111;
    rom_data[2483]=16'b1000100101001111;
    rom_data[2484]=16'b0111010110010010;
    rom_data[2485]=16'b1000100111100110;
    rom_data[2486]=16'b0111010101110101;
    rom_data[2487]=16'b1000101001110001;
    rom_data[2488]=16'b0111010101011000;
    rom_data[2489]=16'b1000101011101110;
    rom_data[2490]=16'b0111010100111010;
    rom_data[2491]=16'b1000101101011100;
    rom_data[2492]=16'b0111010100011101;
    rom_data[2493]=16'b1000101110111011;
    rom_data[2494]=16'b0111010100000000;
    rom_data[2495]=16'b1000110000001010;
    rom_data[2496]=16'b0111010011100011;
    rom_data[2497]=16'b1000110001001001;
    rom_data[2498]=16'b0111010011000110;
    rom_data[2499]=16'b1000110001110111;
    rom_data[2500]=16'b0111010010101010;
    rom_data[2501]=16'b1000110010010100;
    rom_data[2502]=16'b0111010010001101;
    rom_data[2503]=16'b1000110010100000;
    rom_data[2504]=16'b0111010001110001;
    rom_data[2505]=16'b1000110010011010;
    rom_data[2506]=16'b0111010001010101;
    rom_data[2507]=16'b1000110010000011;
    rom_data[2508]=16'b0111010000111001;
    rom_data[2509]=16'b1000110001011010;
    rom_data[2510]=16'b0111010000011110;
    rom_data[2511]=16'b1000110000100000;
    rom_data[2512]=16'b0111010000000011;
    rom_data[2513]=16'b1000101111010110;
    rom_data[2514]=16'b0111001111101000;
    rom_data[2515]=16'b1000101101111011;
    rom_data[2516]=16'b0111001111001110;
    rom_data[2517]=16'b1000101100010000;
    rom_data[2518]=16'b0111001110110011;
    rom_data[2519]=16'b1000101010010111;
    rom_data[2520]=16'b0111001110011010;
    rom_data[2521]=16'b1000101000001111;
    rom_data[2522]=16'b0111001110000000;
    rom_data[2523]=16'b1000100101111001;
    rom_data[2524]=16'b0111001101100111;
    rom_data[2525]=16'b1000100011010110;
    rom_data[2526]=16'b0111001101001110;
    rom_data[2527]=16'b1000100000100111;
    rom_data[2528]=16'b0111001100110101;
    rom_data[2529]=16'b1000011101101101;
    rom_data[2530]=16'b0111001100011101;
    rom_data[2531]=16'b1000011010101000;
    rom_data[2532]=16'b0111001100000100;
    rom_data[2533]=16'b1000010111011001;
    rom_data[2534]=16'b0111001011101100;
    rom_data[2535]=16'b1000010100000000;
    rom_data[2536]=16'b0111001011010101;
    rom_data[2537]=16'b1000010000011110;
    rom_data[2538]=16'b0111001010111101;
    rom_data[2539]=16'b1000001100110101;
    rom_data[2540]=16'b0111001010100110;
    rom_data[2541]=16'b1000001001000011;
    rom_data[2542]=16'b0111001010001111;
    rom_data[2543]=16'b1000000101001011;
    rom_data[2544]=16'b0111001001111000;
    rom_data[2545]=16'b1000000001001100;
    rom_data[2546]=16'b0111001001100010;
    rom_data[2547]=16'b0111111101000111;
    rom_data[2548]=16'b0111001001001011;
    rom_data[2549]=16'b0111111000111100;
    rom_data[2550]=16'b0111001000110101;
    rom_data[2551]=16'b0111110100101100;
    rom_data[2552]=16'b0111001000011111;
    rom_data[2553]=16'b0111110000010111;
    rom_data[2554]=16'b0111001000001001;
    rom_data[2555]=16'b0111101011111110;
    rom_data[2556]=16'b0111000111110011;
    rom_data[2557]=16'b0111100111100000;
    rom_data[2558]=16'b0111000111011110;
    rom_data[2559]=16'b0111100010111110;
    rom_data[2560]=16'b0111000111001000;
    rom_data[2561]=16'b0111011110011001;
    rom_data[2562]=16'b0111000110110011;
    rom_data[2563]=16'b0111011001110001;
    rom_data[2564]=16'b0111000110011101;
    rom_data[2565]=16'b0111010101000101;
    rom_data[2566]=16'b0111000110001000;
    rom_data[2567]=16'b0111010000010111;
    rom_data[2568]=16'b0111000101110011;
    rom_data[2569]=16'b0111001011100110;
    rom_data[2570]=16'b0111000101011110;
    rom_data[2571]=16'b0111000110110011;
    rom_data[2572]=16'b0111000101001001;
    rom_data[2573]=16'b0111000001111101;
    rom_data[2574]=16'b0111000100110100;
    rom_data[2575]=16'b0110111101000101;
    rom_data[2576]=16'b0111000100011111;
    rom_data[2577]=16'b0110111000001100;
    rom_data[2578]=16'b0111000100001011;
    rom_data[2579]=16'b0110110011010001;
    rom_data[2580]=16'b0111000011110110;
    rom_data[2581]=16'b0110101110010100;
    rom_data[2582]=16'b0111000011100001;
    rom_data[2583]=16'b0110101001010110;
    rom_data[2584]=16'b0111000011001100;
    rom_data[2585]=16'b0110100100010111;
    rom_data[2586]=16'b0111000010111000;
    rom_data[2587]=16'b0110011111010111;
    rom_data[2588]=16'b0111000010100011;
    rom_data[2589]=16'b0110011010010101;
    rom_data[2590]=16'b0111000010001110;
    rom_data[2591]=16'b0110010101010011;
    rom_data[2592]=16'b0111000001111010;
    rom_data[2593]=16'b0110010000010001;
    rom_data[2594]=16'b0111000001100101;
    rom_data[2595]=16'b0110001011001101;
    rom_data[2596]=16'b0111000001010000;
    rom_data[2597]=16'b0110000110001010;
    rom_data[2598]=16'b0111000000111100;
    rom_data[2599]=16'b0110000001000110;
    rom_data[2600]=16'b0111000000100111;
    rom_data[2601]=16'b0101111100000010;
    rom_data[2602]=16'b0111000000010010;
    rom_data[2603]=16'b0101110110111110;
    rom_data[2604]=16'b0110111111111101;
    rom_data[2605]=16'b0101110001111001;
    rom_data[2606]=16'b0110111111101000;
    rom_data[2607]=16'b0101101100110110;
    rom_data[2608]=16'b0110111111010011;
    rom_data[2609]=16'b0101100111110010;
    rom_data[2610]=16'b0110111110111110;
    rom_data[2611]=16'b0101100010101111;
    rom_data[2612]=16'b0110111110101001;
    rom_data[2613]=16'b0101011101101100;
    rom_data[2614]=16'b0110111110010100;
    rom_data[2615]=16'b0101011000101010;
    rom_data[2616]=16'b0110111101111111;
    rom_data[2617]=16'b0101010011101001;
    rom_data[2618]=16'b0110111101101001;
    rom_data[2619]=16'b0101001110101000;
    rom_data[2620]=16'b0110111101010100;
    rom_data[2621]=16'b0101001001101001;
    rom_data[2622]=16'b0110111100111110;
    rom_data[2623]=16'b0101000100101011;
    rom_data[2624]=16'b0110111100101000;
    rom_data[2625]=16'b0100111111101110;
    rom_data[2626]=16'b0110111100010010;
    rom_data[2627]=16'b0100111010110011;
    rom_data[2628]=16'b0110111011111100;
    rom_data[2629]=16'b0100110101111001;
    rom_data[2630]=16'b0110111011100110;
    rom_data[2631]=16'b0100110001000001;
    rom_data[2632]=16'b0110111011010000;
    rom_data[2633]=16'b0100101100001011;
    rom_data[2634]=16'b0110111010111001;
    rom_data[2635]=16'b0100100111010111;
    rom_data[2636]=16'b0110111010100010;
    rom_data[2637]=16'b0100100010100110;
    rom_data[2638]=16'b0110111010001011;
    rom_data[2639]=16'b0100011101110111;
    rom_data[2640]=16'b0110111001110100;
    rom_data[2641]=16'b0100011001001010;
    rom_data[2642]=16'b0110111001011101;
    rom_data[2643]=16'b0100010100100001;
    rom_data[2644]=16'b0110111001000101;
    rom_data[2645]=16'b0100001111111010;
    rom_data[2646]=16'b0110111000101101;
    rom_data[2647]=16'b0100001011010111;
    rom_data[2648]=16'b0110111000010101;
    rom_data[2649]=16'b0100000110111000;
    rom_data[2650]=16'b0110110111111100;
    rom_data[2651]=16'b0100000010011101;
    rom_data[2652]=16'b0110110111100100;
    rom_data[2653]=16'b0011111110000101;
    rom_data[2654]=16'b0110110111001010;
    rom_data[2655]=16'b0011111001110011;
    rom_data[2656]=16'b0110110110110001;
    rom_data[2657]=16'b0011110101100101;
    rom_data[2658]=16'b0110110110011000;
    rom_data[2659]=16'b0011110001011100;
    rom_data[2660]=16'b0110110101111110;
    rom_data[2661]=16'b0011101101011001;
    rom_data[2662]=16'b0110110101100011;
    rom_data[2663]=16'b0011101001011100;
    rom_data[2664]=16'b0110110101001001;
    rom_data[2665]=16'b0011100101100101;
    rom_data[2666]=16'b0110110100101110;
    rom_data[2667]=16'b0011100001110101;
    rom_data[2668]=16'b0110110100010011;
    rom_data[2669]=16'b0011011110001101;
    rom_data[2670]=16'b0110110011110111;
    rom_data[2671]=16'b0011011010101100;
    rom_data[2672]=16'b0110110011011011;
    rom_data[2673]=16'b0011010111010100;
    rom_data[2674]=16'b0110110010111111;
    rom_data[2675]=16'b0011010100000101;
    rom_data[2676]=16'b0110110010100011;
    rom_data[2677]=16'b0011010001000000;
    rom_data[2678]=16'b0110110010000111;
    rom_data[2679]=16'b0011001110000101;
    rom_data[2680]=16'b0110110001101010;
    rom_data[2681]=16'b0011001011010101;
    rom_data[2682]=16'b0110110001001101;
    rom_data[2683]=16'b0011001000110001;
    rom_data[2684]=16'b0110110000110000;
    rom_data[2685]=16'b0011000110011010;
    rom_data[2686]=16'b0110110000010011;
    rom_data[2687]=16'b0011000100001111;
    rom_data[2688]=16'b0110101111110110;
    rom_data[2689]=16'b0011000010010010;
    rom_data[2690]=16'b0110101111011000;
    rom_data[2691]=16'b0011000000100100;
    rom_data[2692]=16'b0110101110111011;
    rom_data[2693]=16'b0010111111000101;
    rom_data[2694]=16'b0110101110011110;
    rom_data[2695]=16'b0010111101110110;
    rom_data[2696]=16'b0110101110000001;
    rom_data[2697]=16'b0010111100110111;
    rom_data[2698]=16'b0110101101100100;
    rom_data[2699]=16'b0010111100001001;
    rom_data[2700]=16'b0110101101001000;
    rom_data[2701]=16'b0010111011101100;
    rom_data[2702]=16'b0110101100101011;
    rom_data[2703]=16'b0010111011100000;
    rom_data[2704]=16'b0110101100001111;
    rom_data[2705]=16'b0010111011100110;
    rom_data[2706]=16'b0110101011110011;
    rom_data[2707]=16'b0010111011111101;
    rom_data[2708]=16'b0110101011010111;
    rom_data[2709]=16'b0010111100100110;
    rom_data[2710]=16'b0110101010111100;
    rom_data[2711]=16'b0010111101100000;
    rom_data[2712]=16'b0110101010100001;
    rom_data[2713]=16'b0010111110101010;
    rom_data[2714]=16'b0110101010000110;
    rom_data[2715]=16'b0011000000000101;
    rom_data[2716]=16'b0110101001101011;
    rom_data[2717]=16'b0011000001110000;
    rom_data[2718]=16'b0110101001010001;
    rom_data[2719]=16'b0011000011101001;
    rom_data[2720]=16'b0110101000110111;
    rom_data[2721]=16'b0011000101110001;
    rom_data[2722]=16'b0110101000011110;
    rom_data[2723]=16'b0011001000000111;
    rom_data[2724]=16'b0110101000000101;
    rom_data[2725]=16'b0011001010101010;
    rom_data[2726]=16'b0110100111101100;
    rom_data[2727]=16'b0011001101011001;
    rom_data[2728]=16'b0110100111010011;
    rom_data[2729]=16'b0011010000010011;
    rom_data[2730]=16'b0110100110111010;
    rom_data[2731]=16'b0011010011011000;
    rom_data[2732]=16'b0110100110100010;
    rom_data[2733]=16'b0011010110101000;
    rom_data[2734]=16'b0110100110001010;
    rom_data[2735]=16'b0011011010000000;
    rom_data[2736]=16'b0110100101110011;
    rom_data[2737]=16'b0011011101100010;
    rom_data[2738]=16'b0110100101011011;
    rom_data[2739]=16'b0011100001001100;
    rom_data[2740]=16'b0110100101000100;
    rom_data[2741]=16'b0011100100111101;
    rom_data[2742]=16'b0110100100101101;
    rom_data[2743]=16'b0011101000110101;
    rom_data[2744]=16'b0110100100010110;
    rom_data[2745]=16'b0011101100110100;
    rom_data[2746]=16'b0110100100000000;
    rom_data[2747]=16'b0011110000111001;
    rom_data[2748]=16'b0110100011101001;
    rom_data[2749]=16'b0011110101000100;
    rom_data[2750]=16'b0110100011010011;
    rom_data[2751]=16'b0011111001010100;
    rom_data[2752]=16'b0110100010111101;
    rom_data[2753]=16'b0011111101101001;
    rom_data[2754]=16'b0110100010100111;
    rom_data[2755]=16'b0100000010000011;
    rom_data[2756]=16'b0110100010010001;
    rom_data[2757]=16'b0100000110100000;
    rom_data[2758]=16'b0110100001111100;
    rom_data[2759]=16'b0100001011000010;
    rom_data[2760]=16'b0110100001100110;
    rom_data[2761]=16'b0100001111100111;
    rom_data[2762]=16'b0110100001010001;
    rom_data[2763]=16'b0100010100001111;
    rom_data[2764]=16'b0110100000111011;
    rom_data[2765]=16'b0100011000111011;
    rom_data[2766]=16'b0110100000100110;
    rom_data[2767]=16'b0100011101101001;
    rom_data[2768]=16'b0110100000010001;
    rom_data[2769]=16'b0100100010011010;
    rom_data[2770]=16'b0110011111111100;
    rom_data[2771]=16'b0100100111001110;
    rom_data[2772]=16'b0110011111100111;
    rom_data[2773]=16'b0100101100000011;
    rom_data[2774]=16'b0110011111010010;
    rom_data[2775]=16'b0100110000111011;
    rom_data[2776]=16'b0110011110111101;
    rom_data[2777]=16'b0100110101110100;
    rom_data[2778]=16'b0110011110101001;
    rom_data[2779]=16'b0100111010101111;
    rom_data[2780]=16'b0110011110010100;
    rom_data[2781]=16'b0100111111101100;
    rom_data[2782]=16'b0110011101111111;
    rom_data[2783]=16'b0101000100101010;
    rom_data[2784]=16'b0110011101101010;
    rom_data[2785]=16'b0101001001101001;
    rom_data[2786]=16'b0110011101010110;
    rom_data[2787]=16'b0101001110101010;
    rom_data[2788]=16'b0110011101000001;
    rom_data[2789]=16'b0101010011101011;
    rom_data[2790]=16'b0110011100101100;
    rom_data[2791]=16'b0101011000101101;
    rom_data[2792]=16'b0110011100011000;
    rom_data[2793]=16'b0101011101110000;
    rom_data[2794]=16'b0110011100000011;
    rom_data[2795]=16'b0101100010110011;
    rom_data[2796]=16'b0110011011101110;
    rom_data[2797]=16'b0101100111110110;
    rom_data[2798]=16'b0110011011011010;
    rom_data[2799]=16'b0101101100111010;
    rom_data[2800]=16'b0110011011000101;
    rom_data[2801]=16'b0101110001111110;
    rom_data[2802]=16'b0110011010110000;
    rom_data[2803]=16'b0101110111000011;
    rom_data[2804]=16'b0110011010011011;
    rom_data[2805]=16'b0101111100000111;
    rom_data[2806]=16'b0110011010000110;
    rom_data[2807]=16'b0110000001001011;
    rom_data[2808]=16'b0110011001110001;
    rom_data[2809]=16'b0110000110001110;
    rom_data[2810]=16'b0110011001011100;
    rom_data[2811]=16'b0110001011010010;
    rom_data[2812]=16'b0110011001000111;
    rom_data[2813]=16'b0110010000010100;
    rom_data[2814]=16'b0110011000110010;
    rom_data[2815]=16'b0110010101010110;
    rom_data[2816]=16'b0110011000011101;
    rom_data[2817]=16'b0110011010010111;
    rom_data[2818]=16'b0110011000000111;
    rom_data[2819]=16'b0110011111011000;
    rom_data[2820]=16'b0110010111110010;
    rom_data[2821]=16'b0110100100010111;
    rom_data[2822]=16'b0110010111011100;
    rom_data[2823]=16'b0110101001010101;
    rom_data[2824]=16'b0110010111000110;
    rom_data[2825]=16'b0110101110010010;
    rom_data[2826]=16'b0110010110110000;
    rom_data[2827]=16'b0110110011001101;
    rom_data[2828]=16'b0110010110011010;
    rom_data[2829]=16'b0110111000000111;
    rom_data[2830]=16'b0110010110000100;
    rom_data[2831]=16'b0110111100111111;
    rom_data[2832]=16'b0110010101101110;
    rom_data[2833]=16'b0111000001110101;
    rom_data[2834]=16'b0110010101010111;
    rom_data[2835]=16'b0111000110101001;
    rom_data[2836]=16'b0110010101000000;
    rom_data[2837]=16'b0111001011011010;
    rom_data[2838]=16'b0110010100101001;
    rom_data[2839]=16'b0111010000001001;
    rom_data[2840]=16'b0110010100010010;
    rom_data[2841]=16'b0111010100110110;
    rom_data[2842]=16'b0110010011111011;
    rom_data[2843]=16'b0111011001011111;
    rom_data[2844]=16'b0110010011100011;
    rom_data[2845]=16'b0111011110000110;
    rom_data[2846]=16'b0110010011001011;
    rom_data[2847]=16'b0111100010101001;
    rom_data[2848]=16'b0110010010110011;
    rom_data[2849]=16'b0111100111001000;
    rom_data[2850]=16'b0110010010011010;
    rom_data[2851]=16'b0111101011100100;
    rom_data[2852]=16'b0110010010000001;
    rom_data[2853]=16'b0111101111111011;
    rom_data[2854]=16'b0110010001101000;
    rom_data[2855]=16'b0111110100001110;
    rom_data[2856]=16'b0110010001001111;
    rom_data[2857]=16'b0111111000011100;
    rom_data[2858]=16'b0110010000110101;
    rom_data[2859]=16'b0111111100100100;
    rom_data[2860]=16'b0110010000011100;
    rom_data[2861]=16'b1000000000100111;
    rom_data[2862]=16'b0110010000000001;
    rom_data[2863]=16'b1000000100100100;
    rom_data[2864]=16'b0110001111100111;
    rom_data[2865]=16'b1000001000011011;
    rom_data[2866]=16'b0110001111001100;
    rom_data[2867]=16'b1000001100001011;
    rom_data[2868]=16'b0110001110110001;
    rom_data[2869]=16'b1000001111110011;
    rom_data[2870]=16'b0110001110010101;
    rom_data[2871]=16'b1000010011010100;
    rom_data[2872]=16'b0110001101111001;
    rom_data[2873]=16'b1000010110101100;
    rom_data[2874]=16'b0110001101011101;
    rom_data[2875]=16'b1000011001111011;
    rom_data[2876]=16'b0110001101000001;
    rom_data[2877]=16'b1000011101000000;
    rom_data[2878]=16'b0110001100100101;
    rom_data[2879]=16'b1000011111111011;
    rom_data[2880]=16'b0110001100001000;
    rom_data[2881]=16'b1000100010101011;
    rom_data[2882]=16'b0110001011101011;
    rom_data[2883]=16'b1000100101001111;
    rom_data[2884]=16'b0110001011001110;
    rom_data[2885]=16'b1000100111100111;
    rom_data[2886]=16'b0110001010110001;
    rom_data[2887]=16'b1000101001110001;
    rom_data[2888]=16'b0110001010010100;
    rom_data[2889]=16'b1000101011101110;
    rom_data[2890]=16'b0110001001110110;
    rom_data[2891]=16'b1000101101011100;
    rom_data[2892]=16'b0110001001011001;
    rom_data[2893]=16'b1000101110111011;
    rom_data[2894]=16'b0110001000111100;
    rom_data[2895]=16'b1000110000001010;
    rom_data[2896]=16'b0110001000011111;
    rom_data[2897]=16'b1000110001001001;
    rom_data[2898]=16'b0110001000000010;
    rom_data[2899]=16'b1000110001110111;
    rom_data[2900]=16'b0110000111100110;
    rom_data[2901]=16'b1000110010010100;
    rom_data[2902]=16'b0110000111001001;
    rom_data[2903]=16'b1000110010100000;
    rom_data[2904]=16'b0110000110101101;
    rom_data[2905]=16'b1000110010011010;
    rom_data[2906]=16'b0110000110010001;
    rom_data[2907]=16'b1000110010000011;
    rom_data[2908]=16'b0110000101110101;
    rom_data[2909]=16'b1000110001011010;
    rom_data[2910]=16'b0110000101011010;
    rom_data[2911]=16'b1000110000100000;
    rom_data[2912]=16'b0110000100111111;
    rom_data[2913]=16'b1000101111010101;
    rom_data[2914]=16'b0110000100100100;
    rom_data[2915]=16'b1000101101111011;
    rom_data[2916]=16'b0110000100001001;
    rom_data[2917]=16'b1000101100010000;
    rom_data[2918]=16'b0110000011101111;
    rom_data[2919]=16'b1000101010010111;
    rom_data[2920]=16'b0110000011010101;
    rom_data[2921]=16'b1000101000001111;
    rom_data[2922]=16'b0110000010111100;
    rom_data[2923]=16'b1000100101111001;
    rom_data[2924]=16'b0110000010100011;
    rom_data[2925]=16'b1000100011010110;
    rom_data[2926]=16'b0110000010001010;
    rom_data[2927]=16'b1000100000100111;
    rom_data[2928]=16'b0110000001110001;
    rom_data[2929]=16'b1000011101101101;
    rom_data[2930]=16'b0110000001011000;
    rom_data[2931]=16'b1000011010101000;
    rom_data[2932]=16'b0110000001000000;
    rom_data[2933]=16'b1000010111011000;
    rom_data[2934]=16'b0110000000101000;
    rom_data[2935]=16'b1000010100000000;
    rom_data[2936]=16'b0110000000010001;
    rom_data[2937]=16'b1000010000011110;
    rom_data[2938]=16'b0101111111111001;
    rom_data[2939]=16'b1000001100110100;
    rom_data[2940]=16'b0101111111100010;
    rom_data[2941]=16'b1000001001000011;
    rom_data[2942]=16'b0101111111001011;
    rom_data[2943]=16'b1000000101001011;
    rom_data[2944]=16'b0101111110110100;
    rom_data[2945]=16'b1000000001001100;
    rom_data[2946]=16'b0101111110011110;
    rom_data[2947]=16'b0111111101000111;
    rom_data[2948]=16'b0101111110000111;
    rom_data[2949]=16'b0111111000111100;
    rom_data[2950]=16'b0101111101110001;
    rom_data[2951]=16'b0111110100101100;
    rom_data[2952]=16'b0101111101011011;
    rom_data[2953]=16'b0111110000010111;
    rom_data[2954]=16'b0101111101000101;
    rom_data[2955]=16'b0111101011111101;
    rom_data[2956]=16'b0101111100101111;
    rom_data[2957]=16'b0111100111100000;
    rom_data[2958]=16'b0101111100011010;
    rom_data[2959]=16'b0111100010111110;
    rom_data[2960]=16'b0101111100000100;
    rom_data[2961]=16'b0111011110011001;
    rom_data[2962]=16'b0101111011101111;
    rom_data[2963]=16'b0111011001110001;
    rom_data[2964]=16'b0101111011011001;
    rom_data[2965]=16'b0111010101000101;
    rom_data[2966]=16'b0101111011000100;
    rom_data[2967]=16'b0111010000010111;
    rom_data[2968]=16'b0101111010101111;
    rom_data[2969]=16'b0111001011100110;
    rom_data[2970]=16'b0101111010011010;
    rom_data[2971]=16'b0111000110110010;
    rom_data[2972]=16'b0101111010000101;
    rom_data[2973]=16'b0111000001111101;
    rom_data[2974]=16'b0101111001110000;
    rom_data[2975]=16'b0110111101000101;
    rom_data[2976]=16'b0101111001011011;
    rom_data[2977]=16'b0110111000001100;
    rom_data[2978]=16'b0101111001000110;
    rom_data[2979]=16'b0110110011010000;
    rom_data[2980]=16'b0101111000110010;
    rom_data[2981]=16'b0110101110010100;
    rom_data[2982]=16'b0101111000011101;
    rom_data[2983]=16'b0110101001010110;
    rom_data[2984]=16'b0101111000001000;
    rom_data[2985]=16'b0110100100010110;
    rom_data[2986]=16'b0101110111110100;
    rom_data[2987]=16'b0110011111010110;
    rom_data[2988]=16'b0101110111011111;
    rom_data[2989]=16'b0110011010010101;
    rom_data[2990]=16'b0101110111001010;
    rom_data[2991]=16'b0110010101010011;
    rom_data[2992]=16'b0101110110110110;
    rom_data[2993]=16'b0110010000010000;
    rom_data[2994]=16'b0101110110100001;
    rom_data[2995]=16'b0110001011001101;
    rom_data[2996]=16'b0101110110001100;
    rom_data[2997]=16'b0110000110001001;
    rom_data[2998]=16'b0101110101111000;
    rom_data[2999]=16'b0110000001000110;
    rom_data[3000]=16'b0101110101100011;
    rom_data[3001]=16'b0101111100000001;
    rom_data[3002]=16'b0101110101001110;
    rom_data[3003]=16'b0101110110111101;
    rom_data[3004]=16'b0101110100111001;
    rom_data[3005]=16'b0101110001111001;
    rom_data[3006]=16'b0101110100100100;
    rom_data[3007]=16'b0101101100110101;
    rom_data[3008]=16'b0101110100001111;
    rom_data[3009]=16'b0101100111110010;
    rom_data[3010]=16'b0101110011111010;
    rom_data[3011]=16'b0101100010101110;
    rom_data[3012]=16'b0101110011100101;
    rom_data[3013]=16'b0101011101101100;
    rom_data[3014]=16'b0101110011010000;
    rom_data[3015]=16'b0101011000101010;
    rom_data[3016]=16'b0101110010111011;
    rom_data[3017]=16'b0101010011101000;
    rom_data[3018]=16'b0101110010100101;
    rom_data[3019]=16'b0101001110101000;
    rom_data[3020]=16'b0101110010010000;
    rom_data[3021]=16'b0101001001101001;
    rom_data[3022]=16'b0101110001111010;
    rom_data[3023]=16'b0101000100101011;
    rom_data[3024]=16'b0101110001100100;
    rom_data[3025]=16'b0100111111101110;
    rom_data[3026]=16'b0101110001001110;
    rom_data[3027]=16'b0100111010110011;
    rom_data[3028]=16'b0101110000111000;
    rom_data[3029]=16'b0100110101111001;
    rom_data[3030]=16'b0101110000100010;
    rom_data[3031]=16'b0100110001000001;
    rom_data[3032]=16'b0101110000001100;
    rom_data[3033]=16'b0100101100001011;
    rom_data[3034]=16'b0101101111110101;
    rom_data[3035]=16'b0100100111010111;
    rom_data[3036]=16'b0101101111011110;
    rom_data[3037]=16'b0100100010100101;
    rom_data[3038]=16'b0101101111000111;
    rom_data[3039]=16'b0100011101110110;
    rom_data[3040]=16'b0101101110110000;
    rom_data[3041]=16'b0100011001001010;
    rom_data[3042]=16'b0101101110011000;
    rom_data[3043]=16'b0100010100100000;
    rom_data[3044]=16'b0101101110000001;
    rom_data[3045]=16'b0100001111111010;
    rom_data[3046]=16'b0101101101101001;
    rom_data[3047]=16'b0100001011010111;
    rom_data[3048]=16'b0101101101010001;
    rom_data[3049]=16'b0100000110111000;
    rom_data[3050]=16'b0101101100111000;
    rom_data[3051]=16'b0100000010011100;
    rom_data[3052]=16'b0101101100011111;
    rom_data[3053]=16'b0011111110000101;
    rom_data[3054]=16'b0101101100000110;
    rom_data[3055]=16'b0011111001110010;
    rom_data[3056]=16'b0101101011101101;
    rom_data[3057]=16'b0011110101100100;
    rom_data[3058]=16'b0101101011010011;
    rom_data[3059]=16'b0011110001011100;
    rom_data[3060]=16'b0101101010111001;
    rom_data[3061]=16'b0011101101011000;
    rom_data[3062]=16'b0101101010011111;
    rom_data[3063]=16'b0011101001011011;
    rom_data[3064]=16'b0101101010000101;
    rom_data[3065]=16'b0011100101100101;
    rom_data[3066]=16'b0101101001101010;
    rom_data[3067]=16'b0011100001110101;
    rom_data[3068]=16'b0101101001001111;
    rom_data[3069]=16'b0011011110001100;
    rom_data[3070]=16'b0101101000110011;
    rom_data[3071]=16'b0011011010101100;
    rom_data[3072]=16'b0101101000010111;
    rom_data[3073]=16'b0011010111010100;
    rom_data[3074]=16'b0101100111111011;
    rom_data[3075]=16'b0011010100000101;
    rom_data[3076]=16'b0101100111011111;
    rom_data[3077]=16'b0011010001000000;
    rom_data[3078]=16'b0101100111000010;
    rom_data[3079]=16'b0011001110000101;
    rom_data[3080]=16'b0101100110100110;
    rom_data[3081]=16'b0011001011010101;
    rom_data[3082]=16'b0101100110001001;
    rom_data[3083]=16'b0011001000110001;
    rom_data[3084]=16'b0101100101101100;
    rom_data[3085]=16'b0011000110011001;
    rom_data[3086]=16'b0101100101001111;
    rom_data[3087]=16'b0011000100001111;
    rom_data[3088]=16'b0101100100110001;
    rom_data[3089]=16'b0011000010010010;
    rom_data[3090]=16'b0101100100010100;
    rom_data[3091]=16'b0011000000100100;
    rom_data[3092]=16'b0101100011110111;
    rom_data[3093]=16'b0010111111000101;
    rom_data[3094]=16'b0101100011011010;
    rom_data[3095]=16'b0010111101110110;
    rom_data[3096]=16'b0101100010111101;
    rom_data[3097]=16'b0010111100110111;
    rom_data[3098]=16'b0101100010100000;
    rom_data[3099]=16'b0010111100001001;
    rom_data[3100]=16'b0101100010000011;
    rom_data[3101]=16'b0010111011101100;
    rom_data[3102]=16'b0101100001100111;
    rom_data[3103]=16'b0010111011100000;
    rom_data[3104]=16'b0101100001001011;
    rom_data[3105]=16'b0010111011100110;
    rom_data[3106]=16'b0101100000101111;
    rom_data[3107]=16'b0010111011111101;
    rom_data[3108]=16'b0101100000010011;
    rom_data[3109]=16'b0010111100100110;
    rom_data[3110]=16'b0101011111111000;
    rom_data[3111]=16'b0010111101100000;
    rom_data[3112]=16'b0101011111011101;
    rom_data[3113]=16'b0010111110101011;
    rom_data[3114]=16'b0101011111000010;
    rom_data[3115]=16'b0011000000000101;
    rom_data[3116]=16'b0101011110100111;
    rom_data[3117]=16'b0011000001110000;
    rom_data[3118]=16'b0101011110001101;
    rom_data[3119]=16'b0011000011101010;
    rom_data[3120]=16'b0101011101110011;
    rom_data[3121]=16'b0011000101110010;
    rom_data[3122]=16'b0101011101011010;
    rom_data[3123]=16'b0011001000000111;
    rom_data[3124]=16'b0101011101000000;
    rom_data[3125]=16'b0011001010101010;
    rom_data[3126]=16'b0101011100100111;
    rom_data[3127]=16'b0011001101011001;
    rom_data[3128]=16'b0101011100001111;
    rom_data[3129]=16'b0011010000010011;
    rom_data[3130]=16'b0101011011110110;
    rom_data[3131]=16'b0011010011011001;
    rom_data[3132]=16'b0101011011011110;
    rom_data[3133]=16'b0011010110101000;
    rom_data[3134]=16'b0101011011000110;
    rom_data[3135]=16'b0011011010000001;
    rom_data[3136]=16'b0101011010101111;
    rom_data[3137]=16'b0011011101100010;
    rom_data[3138]=16'b0101011010010111;
    rom_data[3139]=16'b0011100001001100;
    rom_data[3140]=16'b0101011010000000;
    rom_data[3141]=16'b0011100100111101;
    rom_data[3142]=16'b0101011001101001;
    rom_data[3143]=16'b0011101000110110;
    rom_data[3144]=16'b0101011001010010;
    rom_data[3145]=16'b0011101100110101;
    rom_data[3146]=16'b0101011000111100;
    rom_data[3147]=16'b0011110000111010;
    rom_data[3148]=16'b0101011000100101;
    rom_data[3149]=16'b0011110101000100;
    rom_data[3150]=16'b0101011000001111;
    rom_data[3151]=16'b0011111001010100;
    rom_data[3152]=16'b0101010111111001;
    rom_data[3153]=16'b0011111101101001;
    rom_data[3154]=16'b0101010111100011;
    rom_data[3155]=16'b0100000010000011;
    rom_data[3156]=16'b0101010111001101;
    rom_data[3157]=16'b0100000110100001;
    rom_data[3158]=16'b0101010110110111;
    rom_data[3159]=16'b0100001011000010;
    rom_data[3160]=16'b0101010110100010;
    rom_data[3161]=16'b0100001111100111;
    rom_data[3162]=16'b0101010110001101;
    rom_data[3163]=16'b0100010100010000;
    rom_data[3164]=16'b0101010101110111;
    rom_data[3165]=16'b0100011000111011;
    rom_data[3166]=16'b0101010101100010;
    rom_data[3167]=16'b0100011101101010;
    rom_data[3168]=16'b0101010101001101;
    rom_data[3169]=16'b0100100010011011;
    rom_data[3170]=16'b0101010100111000;
    rom_data[3171]=16'b0100100111001110;
    rom_data[3172]=16'b0101010100100011;
    rom_data[3173]=16'b0100101100000100;
    rom_data[3174]=16'b0101010100001110;
    rom_data[3175]=16'b0100110000111011;
    rom_data[3176]=16'b0101010011111001;
    rom_data[3177]=16'b0100110101110101;
    rom_data[3178]=16'b0101010011100100;
    rom_data[3179]=16'b0100111010110000;
    rom_data[3180]=16'b0101010011010000;
    rom_data[3181]=16'b0100111111101100;
    rom_data[3182]=16'b0101010010111011;
    rom_data[3183]=16'b0101000100101010;
    rom_data[3184]=16'b0101010010100110;
    rom_data[3185]=16'b0101001001101010;
    rom_data[3186]=16'b0101010010010010;
    rom_data[3187]=16'b0101001110101010;
    rom_data[3188]=16'b0101010001111101;
    rom_data[3189]=16'b0101010011101011;
    rom_data[3190]=16'b0101010001101000;
    rom_data[3191]=16'b0101011000101101;
    rom_data[3192]=16'b0101010001010100;
    rom_data[3193]=16'b0101011101110000;
    rom_data[3194]=16'b0101010000111111;
    rom_data[3195]=16'b0101100010110011;
    rom_data[3196]=16'b0101010000101010;
    rom_data[3197]=16'b0101100111110111;
    rom_data[3198]=16'b0101010000010110;
    rom_data[3199]=16'b0101101100111011;
    rom_data[3200]=16'b0101010000000001;
    rom_data[3201]=16'b0101110001111111;
    rom_data[3202]=16'b0101001111101100;
    rom_data[3203]=16'b0101110111000011;
    rom_data[3204]=16'b0101001111010111;
    rom_data[3205]=16'b0101111100000111;
    rom_data[3206]=16'b0101001111000010;
    rom_data[3207]=16'b0110000001001011;
    rom_data[3208]=16'b0101001110101101;
    rom_data[3209]=16'b0110000110001111;
    rom_data[3210]=16'b0101001110011000;
    rom_data[3211]=16'b0110001011010010;
    rom_data[3212]=16'b0101001110000011;
    rom_data[3213]=16'b0110010000010101;
    rom_data[3214]=16'b0101001101101110;
    rom_data[3215]=16'b0110010101010111;
    rom_data[3216]=16'b0101001101011001;
    rom_data[3217]=16'b0110011010011000;
    rom_data[3218]=16'b0101001101000011;
    rom_data[3219]=16'b0110011111011000;
    rom_data[3220]=16'b0101001100101110;
    rom_data[3221]=16'b0110100100010111;
    rom_data[3222]=16'b0101001100011000;
    rom_data[3223]=16'b0110101001010110;
    rom_data[3224]=16'b0101001100000010;
    rom_data[3225]=16'b0110101110010010;
    rom_data[3226]=16'b0101001011101100;
    rom_data[3227]=16'b0110110011001110;
    rom_data[3228]=16'b0101001011010110;
    rom_data[3229]=16'b0110111000000111;
    rom_data[3230]=16'b0101001011000000;
    rom_data[3231]=16'b0110111100111111;
    rom_data[3232]=16'b0101001010101010;
    rom_data[3233]=16'b0111000001110101;
    rom_data[3234]=16'b0101001010010011;
    rom_data[3235]=16'b0111000110101001;
    rom_data[3236]=16'b0101001001111100;
    rom_data[3237]=16'b0111001011011011;
    rom_data[3238]=16'b0101001001100101;
    rom_data[3239]=16'b0111010000001010;
    rom_data[3240]=16'b0101001001001110;
    rom_data[3241]=16'b0111010100110110;
    rom_data[3242]=16'b0101001000110110;
    rom_data[3243]=16'b0111011001100000;
    rom_data[3244]=16'b0101001000011111;
    rom_data[3245]=16'b0111011110000110;
    rom_data[3246]=16'b0101001000000111;
    rom_data[3247]=16'b0111100010101001;
    rom_data[3248]=16'b0101000111101111;
    rom_data[3249]=16'b0111100111001000;
    rom_data[3250]=16'b0101000111010110;
    rom_data[3251]=16'b0111101011100100;
    rom_data[3252]=16'b0101000110111101;
    rom_data[3253]=16'b0111101111111011;
    rom_data[3254]=16'b0101000110100100;
    rom_data[3255]=16'b0111110100001110;
    rom_data[3256]=16'b0101000110001011;
    rom_data[3257]=16'b0111111000011100;
    rom_data[3258]=16'b0101000101110001;
    rom_data[3259]=16'b0111111100100101;
    rom_data[3260]=16'b0101000101010111;
    rom_data[3261]=16'b1000000000101000;
    rom_data[3262]=16'b0101000100111101;
    rom_data[3263]=16'b1000000100100101;
    rom_data[3264]=16'b0101000100100011;
    rom_data[3265]=16'b1000001000011011;
    rom_data[3266]=16'b0101000100001000;
    rom_data[3267]=16'b1000001100001011;
    rom_data[3268]=16'b0101000011101101;
    rom_data[3269]=16'b1000001111110100;
    rom_data[3270]=16'b0101000011010001;
    rom_data[3271]=16'b1000010011010100;
    rom_data[3272]=16'b0101000010110101;
    rom_data[3273]=16'b1000010110101100;
    rom_data[3274]=16'b0101000010011001;
    rom_data[3275]=16'b1000011001111011;
    rom_data[3276]=16'b0101000001111101;
    rom_data[3277]=16'b1000011101000000;
    rom_data[3278]=16'b0101000001100000;
    rom_data[3279]=16'b1000011111111011;
    rom_data[3280]=16'b0101000001000100;
    rom_data[3281]=16'b1000100010101011;
    rom_data[3282]=16'b0101000000100111;
    rom_data[3283]=16'b1000100101001111;
    rom_data[3284]=16'b0101000000001010;
    rom_data[3285]=16'b1000100111100111;
    rom_data[3286]=16'b0100111111101101;
    rom_data[3287]=16'b1000101001110001;
    rom_data[3288]=16'b0100111111001111;
    rom_data[3289]=16'b1000101011101110;
    rom_data[3290]=16'b0100111110110010;
    rom_data[3291]=16'b1000101101011100;
    rom_data[3292]=16'b0100111110010101;
    rom_data[3293]=16'b1000101110111011;
    rom_data[3294]=16'b0100111101111000;
    rom_data[3295]=16'b1000110000001010;
    rom_data[3296]=16'b0100111101011011;
    rom_data[3297]=16'b1000110001001001;
    rom_data[3298]=16'b0100111100111110;
    rom_data[3299]=16'b1000110001110111;
    rom_data[3300]=16'b0100111100100001;
    rom_data[3301]=16'b1000110010010100;
    rom_data[3302]=16'b0100111100000101;
    rom_data[3303]=16'b1000110010100000;
    rom_data[3304]=16'b0100111011101001;
    rom_data[3305]=16'b1000110010011010;
    rom_data[3306]=16'b0100111011001101;
    rom_data[3307]=16'b1000110010000011;
    rom_data[3308]=16'b0100111010110001;
    rom_data[3309]=16'b1000110001011010;
    rom_data[3310]=16'b0100111010010110;
    rom_data[3311]=16'b1000110000100000;
    rom_data[3312]=16'b0100111001111011;
    rom_data[3313]=16'b1000101111010101;
    rom_data[3314]=16'b0100111001100000;
    rom_data[3315]=16'b1000101101111011;
    rom_data[3316]=16'b0100111001000101;
    rom_data[3317]=16'b1000101100010000;
    rom_data[3318]=16'b0100111000101011;
    rom_data[3319]=16'b1000101010010110;
    rom_data[3320]=16'b0100111000010001;
    rom_data[3321]=16'b1000101000001110;
    rom_data[3322]=16'b0100110111111000;
    rom_data[3323]=16'b1000100101111001;
    rom_data[3324]=16'b0100110111011110;
    rom_data[3325]=16'b1000100011010110;
    rom_data[3326]=16'b0100110111000101;
    rom_data[3327]=16'b1000100000100111;
    rom_data[3328]=16'b0100110110101101;
    rom_data[3329]=16'b1000011101101101;
    rom_data[3330]=16'b0100110110010100;
    rom_data[3331]=16'b1000011010100111;
    rom_data[3332]=16'b0100110101111100;
    rom_data[3333]=16'b1000010111011000;
    rom_data[3334]=16'b0100110101100100;
    rom_data[3335]=16'b1000010011111111;
    rom_data[3336]=16'b0100110101001101;
    rom_data[3337]=16'b1000010000011110;
    rom_data[3338]=16'b0100110100110101;
    rom_data[3339]=16'b1000001100110100;
    rom_data[3340]=16'b0100110100011110;
    rom_data[3341]=16'b1000001001000011;
    rom_data[3342]=16'b0100110100000111;
    rom_data[3343]=16'b1000000101001010;
    rom_data[3344]=16'b0100110011110000;
    rom_data[3345]=16'b1000000001001011;
    rom_data[3346]=16'b0100110011011010;
    rom_data[3347]=16'b0111111101000110;
    rom_data[3348]=16'b0100110011000011;
    rom_data[3349]=16'b0111111000111011;
    rom_data[3350]=16'b0100110010101101;
    rom_data[3351]=16'b0111110100101011;
    rom_data[3352]=16'b0100110010010111;
    rom_data[3353]=16'b0111110000010110;
    rom_data[3354]=16'b0100110010000001;
    rom_data[3355]=16'b0111101011111101;
    rom_data[3356]=16'b0100110001101011;
    rom_data[3357]=16'b0111100111011111;
    rom_data[3358]=16'b0100110001010101;
    rom_data[3359]=16'b0111100010111110;
    rom_data[3360]=16'b0100110001000000;
    rom_data[3361]=16'b0111011110011001;
    rom_data[3362]=16'b0100110000101010;
    rom_data[3363]=16'b0111011001110000;
    rom_data[3364]=16'b0100110000010101;
    rom_data[3365]=16'b0111010101000101;
    rom_data[3366]=16'b0100110000000000;
    rom_data[3367]=16'b0111010000010110;
    rom_data[3368]=16'b0100101111101011;
    rom_data[3369]=16'b0111001011100101;
    rom_data[3370]=16'b0100101111010110;
    rom_data[3371]=16'b0111000110110010;
    rom_data[3372]=16'b0100101111000001;
    rom_data[3373]=16'b0111000001111100;
    rom_data[3374]=16'b0100101110101100;
    rom_data[3375]=16'b0110111101000101;
    rom_data[3376]=16'b0100101110010111;
    rom_data[3377]=16'b0110111000001011;
    rom_data[3378]=16'b0100101110000010;
    rom_data[3379]=16'b0110110011010000;
    rom_data[3380]=16'b0100101101101110;
    rom_data[3381]=16'b0110101110010011;
    rom_data[3382]=16'b0100101101011001;
    rom_data[3383]=16'b0110101001010101;
    rom_data[3384]=16'b0100101101000100;
    rom_data[3385]=16'b0110100100010110;
    rom_data[3386]=16'b0100101100110000;
    rom_data[3387]=16'b0110011111010110;
    rom_data[3388]=16'b0100101100011011;
    rom_data[3389]=16'b0110011010010101;
    rom_data[3390]=16'b0100101100000110;
    rom_data[3391]=16'b0110010101010011;
    rom_data[3392]=16'b0100101011110010;
    rom_data[3393]=16'b0110010000010000;
    rom_data[3394]=16'b0100101011011101;
    rom_data[3395]=16'b0110001011001101;
    rom_data[3396]=16'b0100101011001000;
    rom_data[3397]=16'b0110000110001001;
    rom_data[3398]=16'b0100101010110011;
    rom_data[3399]=16'b0110000001000101;
    rom_data[3400]=16'b0100101010011111;
    rom_data[3401]=16'b0101111100000001;
    rom_data[3402]=16'b0100101010001010;
    rom_data[3403]=16'b0101110110111101;
    rom_data[3404]=16'b0100101001110101;
    rom_data[3405]=16'b0101110001111001;
    rom_data[3406]=16'b0100101001100000;
    rom_data[3407]=16'b0101101100110101;
    rom_data[3408]=16'b0100101001001011;
    rom_data[3409]=16'b0101100111110001;
    rom_data[3410]=16'b0100101000110110;
    rom_data[3411]=16'b0101100010101110;
    rom_data[3412]=16'b0100101000100001;
    rom_data[3413]=16'b0101011101101011;
    rom_data[3414]=16'b0100101000001100;
    rom_data[3415]=16'b0101011000101001;
    rom_data[3416]=16'b0100100111110111;
    rom_data[3417]=16'b0101010011101000;
    rom_data[3418]=16'b0100100111100001;
    rom_data[3419]=16'b0101001110101000;
    rom_data[3420]=16'b0100100111001100;
    rom_data[3421]=16'b0101001001101000;
    rom_data[3422]=16'b0100100110110110;
    rom_data[3423]=16'b0101000100101010;
    rom_data[3424]=16'b0100100110100000;
    rom_data[3425]=16'b0100111111101110;
    rom_data[3426]=16'b0100100110001010;
    rom_data[3427]=16'b0100111010110010;
    rom_data[3428]=16'b0100100101110100;
    rom_data[3429]=16'b0100110101111000;
    rom_data[3430]=16'b0100100101011110;
    rom_data[3431]=16'b0100110001000001;
    rom_data[3432]=16'b0100100101000111;
    rom_data[3433]=16'b0100101100001011;
    rom_data[3434]=16'b0100100100110001;
    rom_data[3435]=16'b0100100111010111;
    rom_data[3436]=16'b0100100100011010;
    rom_data[3437]=16'b0100100010100101;
    rom_data[3438]=16'b0100100100000011;
    rom_data[3439]=16'b0100011101110110;
    rom_data[3440]=16'b0100100011101100;
    rom_data[3441]=16'b0100011001001010;
    rom_data[3442]=16'b0100100011010100;
    rom_data[3443]=16'b0100010100100000;
    rom_data[3444]=16'b0100100010111101;
    rom_data[3445]=16'b0100001111111010;
    rom_data[3446]=16'b0100100010100101;
    rom_data[3447]=16'b0100001011010111;
    rom_data[3448]=16'b0100100010001100;
    rom_data[3449]=16'b0100000110110111;
    rom_data[3450]=16'b0100100001110100;
    rom_data[3451]=16'b0100000010011100;
    rom_data[3452]=16'b0100100001011011;
    rom_data[3453]=16'b0011111110000101;
    rom_data[3454]=16'b0100100001000010;
    rom_data[3455]=16'b0011111001110010;
    rom_data[3456]=16'b0100100000101001;
    rom_data[3457]=16'b0011110101100100;
    rom_data[3458]=16'b0100100000001111;
    rom_data[3459]=16'b0011110001011011;
    rom_data[3460]=16'b0100011111110101;
    rom_data[3461]=16'b0011101101011000;
    rom_data[3462]=16'b0100011111011011;
    rom_data[3463]=16'b0011101001011011;
    rom_data[3464]=16'b0100011111000001;
    rom_data[3465]=16'b0011100101100100;
    rom_data[3466]=16'b0100011110100110;
    rom_data[3467]=16'b0011100001110101;
    rom_data[3468]=16'b0100011110001010;
    rom_data[3469]=16'b0011011110001100;
    rom_data[3470]=16'b0100011101101111;
    rom_data[3471]=16'b0011011010101100;
    rom_data[3472]=16'b0100011101010011;
    rom_data[3473]=16'b0011010111010100;
    rom_data[3474]=16'b0100011100110111;
    rom_data[3475]=16'b0011010100000101;
    rom_data[3476]=16'b0100011100011011;
    rom_data[3477]=16'b0011010001000000;
    rom_data[3478]=16'b0100011011111110;
    rom_data[3479]=16'b0011001110000101;
    rom_data[3480]=16'b0100011011100010;
    rom_data[3481]=16'b0011001011010101;
    rom_data[3482]=16'b0100011011000101;
    rom_data[3483]=16'b0011001000110001;
    rom_data[3484]=16'b0100011010101000;
    rom_data[3485]=16'b0011000110011001;
    rom_data[3486]=16'b0100011010001011;
    rom_data[3487]=16'b0011000100001111;
    rom_data[3488]=16'b0100011001101101;
    rom_data[3489]=16'b0011000010010010;
    rom_data[3490]=16'b0100011001010000;
    rom_data[3491]=16'b0011000000100100;
    rom_data[3492]=16'b0100011000110011;
    rom_data[3493]=16'b0010111111000101;
    rom_data[3494]=16'b0100011000010110;
    rom_data[3495]=16'b0010111101110110;
    rom_data[3496]=16'b0100010111111001;
    rom_data[3497]=16'b0010111100110111;
    rom_data[3498]=16'b0100010111011100;
    rom_data[3499]=16'b0010111100001001;
    rom_data[3500]=16'b0100010110111111;
    rom_data[3501]=16'b0010111011101100;
    rom_data[3502]=16'b0100010110100011;
    rom_data[3503]=16'b0010111011100000;
    rom_data[3504]=16'b0100010110000111;
    rom_data[3505]=16'b0010111011100110;
    rom_data[3506]=16'b0100010101101011;
    rom_data[3507]=16'b0010111011111110;
    rom_data[3508]=16'b0100010101001111;
    rom_data[3509]=16'b0010111100100110;
    rom_data[3510]=16'b0100010100110100;
    rom_data[3511]=16'b0010111101100000;
    rom_data[3512]=16'b0100010100011000;
    rom_data[3513]=16'b0010111110101011;
    rom_data[3514]=16'b0100010011111110;
    rom_data[3515]=16'b0011000000000101;
    rom_data[3516]=16'b0100010011100011;
    rom_data[3517]=16'b0011000001110000;
    rom_data[3518]=16'b0100010011001001;
    rom_data[3519]=16'b0011000011101010;
    rom_data[3520]=16'b0100010010101111;
    rom_data[3521]=16'b0011000101110010;
    rom_data[3522]=16'b0100010010010110;
    rom_data[3523]=16'b0011001000000111;
    rom_data[3524]=16'b0100010001111100;
    rom_data[3525]=16'b0011001010101010;
    rom_data[3526]=16'b0100010001100011;
    rom_data[3527]=16'b0011001101011001;
    rom_data[3528]=16'b0100010001001011;
    rom_data[3529]=16'b0011010000010100;
    rom_data[3530]=16'b0100010000110010;
    rom_data[3531]=16'b0011010011011001;
    rom_data[3532]=16'b0100010000011010;
    rom_data[3533]=16'b0011010110101000;
    rom_data[3534]=16'b0100010000000010;
    rom_data[3535]=16'b0011011010000001;
    rom_data[3536]=16'b0100001111101010;
    rom_data[3537]=16'b0011011101100010;
    rom_data[3538]=16'b0100001111010011;
    rom_data[3539]=16'b0011100001001100;
    rom_data[3540]=16'b0100001110111100;
    rom_data[3541]=16'b0011100100111101;
    rom_data[3542]=16'b0100001110100101;
    rom_data[3543]=16'b0011101000110110;
    rom_data[3544]=16'b0100001110001110;
    rom_data[3545]=16'b0011101100110101;
    rom_data[3546]=16'b0100001101110111;
    rom_data[3547]=16'b0011110000111010;
    rom_data[3548]=16'b0100001101100001;
    rom_data[3549]=16'b0011110101000101;
    rom_data[3550]=16'b0100001101001011;
    rom_data[3551]=16'b0011111001010101;
    rom_data[3552]=16'b0100001100110101;
    rom_data[3553]=16'b0011111101101010;
    rom_data[3554]=16'b0100001100011111;
    rom_data[3555]=16'b0100000010000011;
    rom_data[3556]=16'b0100001100001001;
    rom_data[3557]=16'b0100000110100001;
    rom_data[3558]=16'b0100001011110011;
    rom_data[3559]=16'b0100001011000010;
    rom_data[3560]=16'b0100001011011110;
    rom_data[3561]=16'b0100001111101000;
    rom_data[3562]=16'b0100001011001000;
    rom_data[3563]=16'b0100010100010000;
    rom_data[3564]=16'b0100001010110011;
    rom_data[3565]=16'b0100011000111100;
    rom_data[3566]=16'b0100001010011110;
    rom_data[3567]=16'b0100011101101010;
    rom_data[3568]=16'b0100001010001001;
    rom_data[3569]=16'b0100100010011011;
    rom_data[3570]=16'b0100001001110100;
    rom_data[3571]=16'b0100100111001110;
    rom_data[3572]=16'b0100001001011111;
    rom_data[3573]=16'b0100101100000100;
    rom_data[3574]=16'b0100001001001010;
    rom_data[3575]=16'b0100110000111100;
    rom_data[3576]=16'b0100001000110101;
    rom_data[3577]=16'b0100110101110101;
    rom_data[3578]=16'b0100001000100000;
    rom_data[3579]=16'b0100111010110000;
    rom_data[3580]=16'b0100001000001100;
    rom_data[3581]=16'b0100111111101101;
    rom_data[3582]=16'b0100000111110111;
    rom_data[3583]=16'b0101000100101011;
    rom_data[3584]=16'b0100000111100010;
    rom_data[3585]=16'b0101001001101010;
    rom_data[3586]=16'b0100000111001101;
    rom_data[3587]=16'b0101001110101010;
    rom_data[3588]=16'b0100000110111001;
    rom_data[3589]=16'b0101010011101100;
    rom_data[3590]=16'b0100000110100100;
    rom_data[3591]=16'b0101011000101110;
    rom_data[3592]=16'b0100000110001111;
    rom_data[3593]=16'b0101011101110000;
    rom_data[3594]=16'b0100000101111011;
    rom_data[3595]=16'b0101100010110011;
    rom_data[3596]=16'b0100000101100110;
    rom_data[3597]=16'b0101100111110111;
    rom_data[3598]=16'b0100000101010001;
    rom_data[3599]=16'b0101101100111011;
    rom_data[3600]=16'b0100000100111101;
    rom_data[3601]=16'b0101110001111111;
    rom_data[3602]=16'b0100000100101000;
    rom_data[3603]=16'b0101110111000011;
    rom_data[3604]=16'b0100000100010011;
    rom_data[3605]=16'b0101111100000111;
    rom_data[3606]=16'b0100000011111110;
    rom_data[3607]=16'b0110000001001011;
    rom_data[3608]=16'b0100000011101001;
    rom_data[3609]=16'b0110000110001111;
    rom_data[3610]=16'b0100000011010100;
    rom_data[3611]=16'b0110001011010010;
    rom_data[3612]=16'b0100000010111111;
    rom_data[3613]=16'b0110010000010101;
    rom_data[3614]=16'b0100000010101010;
    rom_data[3615]=16'b0110010101010111;
    rom_data[3616]=16'b0100000010010100;
    rom_data[3617]=16'b0110011010011000;
    rom_data[3618]=16'b0100000001111111;
    rom_data[3619]=16'b0110011111011001;
    rom_data[3620]=16'b0100000001101010;
    rom_data[3621]=16'b0110100100011000;
    rom_data[3622]=16'b0100000001010100;
    rom_data[3623]=16'b0110101001010110;
    rom_data[3624]=16'b0100000000111110;
    rom_data[3625]=16'b0110101110010011;
    rom_data[3626]=16'b0100000000101000;
    rom_data[3627]=16'b0110110011001110;
    rom_data[3628]=16'b0100000000010010;
    rom_data[3629]=16'b0110111000001000;
    rom_data[3630]=16'b0011111111111100;
    rom_data[3631]=16'b0110111101000000;
    rom_data[3632]=16'b0011111111100101;
    rom_data[3633]=16'b0111000001110110;
    rom_data[3634]=16'b0011111111001111;
    rom_data[3635]=16'b0111000110101001;
    rom_data[3636]=16'b0011111110111000;
    rom_data[3637]=16'b0111001011011011;
    rom_data[3638]=16'b0011111110100001;
    rom_data[3639]=16'b0111010000001010;
    rom_data[3640]=16'b0011111110001010;
    rom_data[3641]=16'b0111010100110111;
    rom_data[3642]=16'b0011111101110010;
    rom_data[3643]=16'b0111011001100000;
    rom_data[3644]=16'b0011111101011011;
    rom_data[3645]=16'b0111011110000110;
    rom_data[3646]=16'b0011111101000011;
    rom_data[3647]=16'b0111100010101001;
    rom_data[3648]=16'b0011111100101010;
    rom_data[3649]=16'b0111100111001001;
    rom_data[3650]=16'b0011111100010010;
    rom_data[3651]=16'b0111101011100100;
    rom_data[3652]=16'b0011111011111001;
    rom_data[3653]=16'b0111101111111011;
    rom_data[3654]=16'b0011111011100000;
    rom_data[3655]=16'b0111110100001110;
    rom_data[3656]=16'b0011111011000111;
    rom_data[3657]=16'b0111111000011100;
    rom_data[3658]=16'b0011111010101101;
    rom_data[3659]=16'b0111111100100101;
    rom_data[3660]=16'b0011111010010011;
    rom_data[3661]=16'b1000000000101000;
    rom_data[3662]=16'b0011111001111001;
    rom_data[3663]=16'b1000000100100101;
    rom_data[3664]=16'b0011111001011110;
    rom_data[3665]=16'b1000001000011100;
    rom_data[3666]=16'b0011111001000100;
    rom_data[3667]=16'b1000001100001100;
    rom_data[3668]=16'b0011111000101000;
    rom_data[3669]=16'b1000001111110100;
    rom_data[3670]=16'b0011111000001101;
    rom_data[3671]=16'b1000010011010100;
    rom_data[3672]=16'b0011110111110001;
    rom_data[3673]=16'b1000010110101100;
    rom_data[3674]=16'b0011110111010101;
    rom_data[3675]=16'b1000011001111011;
    rom_data[3676]=16'b0011110110111001;
    rom_data[3677]=16'b1000011101000000;
    rom_data[3678]=16'b0011110110011100;
    rom_data[3679]=16'b1000011111111011;
    rom_data[3680]=16'b0011110110000000;
    rom_data[3681]=16'b1000100010101011;
    rom_data[3682]=16'b0011110101100011;
    rom_data[3683]=16'b1000100101001111;
    rom_data[3684]=16'b0011110101000110;
    rom_data[3685]=16'b1000100111100111;
    rom_data[3686]=16'b0011110100101000;
    rom_data[3687]=16'b1000101001110001;
    rom_data[3688]=16'b0011110100001011;
    rom_data[3689]=16'b1000101011101110;
    rom_data[3690]=16'b0011110011101110;
    rom_data[3691]=16'b1000101101011100;
    rom_data[3692]=16'b0011110011010001;
    rom_data[3693]=16'b1000101110111011;
    rom_data[3694]=16'b0011110010110100;
    rom_data[3695]=16'b1000110000001010;
    rom_data[3696]=16'b0011110010010111;
    rom_data[3697]=16'b1000110001001001;
    rom_data[3698]=16'b0011110001111010;
    rom_data[3699]=16'b1000110001110111;
    rom_data[3700]=16'b0011110001011101;
    rom_data[3701]=16'b1000110010010100;
    rom_data[3702]=16'b0011110001000001;
    rom_data[3703]=16'b1000110010100000;
    rom_data[3704]=16'b0011110000100101;
    rom_data[3705]=16'b1000110010011010;
    rom_data[3706]=16'b0011110000001001;
    rom_data[3707]=16'b1000110010000010;
    rom_data[3708]=16'b0011101111101101;
    rom_data[3709]=16'b1000110001011010;
    rom_data[3710]=16'b0011101111010010;
    rom_data[3711]=16'b1000110000100000;
    rom_data[3712]=16'b0011101110110110;
    rom_data[3713]=16'b1000101111010101;
    rom_data[3714]=16'b0011101110011100;
    rom_data[3715]=16'b1000101101111010;
    rom_data[3716]=16'b0011101110000001;
    rom_data[3717]=16'b1000101100010000;
    rom_data[3718]=16'b0011101101100111;
    rom_data[3719]=16'b1000101010010110;
    rom_data[3720]=16'b0011101101001101;
    rom_data[3721]=16'b1000101000001110;
    rom_data[3722]=16'b0011101100110100;
    rom_data[3723]=16'b1000100101111000;
    rom_data[3724]=16'b0011101100011010;
    rom_data[3725]=16'b1000100011010110;
    rom_data[3726]=16'b0011101100000001;
    rom_data[3727]=16'b1000100000100111;
    rom_data[3728]=16'b0011101011101001;
    rom_data[3729]=16'b1000011101101100;
    rom_data[3730]=16'b0011101011010000;
    rom_data[3731]=16'b1000011010100111;
    rom_data[3732]=16'b0011101010111000;
    rom_data[3733]=16'b1000010111011000;
    rom_data[3734]=16'b0011101010100000;
    rom_data[3735]=16'b1000010011111111;
    rom_data[3736]=16'b0011101010001000;
    rom_data[3737]=16'b1000010000011110;
    rom_data[3738]=16'b0011101001110001;
    rom_data[3739]=16'b1000001100110100;
    rom_data[3740]=16'b0011101001011010;
    rom_data[3741]=16'b1000001001000010;
    rom_data[3742]=16'b0011101001000011;
    rom_data[3743]=16'b1000000101001010;
    rom_data[3744]=16'b0011101000101100;
    rom_data[3745]=16'b1000000001001011;
    rom_data[3746]=16'b0011101000010101;
    rom_data[3747]=16'b0111111101000110;
    rom_data[3748]=16'b0011100111111111;
    rom_data[3749]=16'b0111111000111011;
    rom_data[3750]=16'b0011100111101001;
    rom_data[3751]=16'b0111110100101011;
    rom_data[3752]=16'b0011100111010011;
    rom_data[3753]=16'b0111110000010110;
    rom_data[3754]=16'b0011100110111101;
    rom_data[3755]=16'b0111101011111101;
    rom_data[3756]=16'b0011100110100111;
    rom_data[3757]=16'b0111100111011111;
    rom_data[3758]=16'b0011100110010001;
    rom_data[3759]=16'b0111100010111101;
    rom_data[3760]=16'b0011100101111100;
    rom_data[3761]=16'b0111011110011000;
    rom_data[3762]=16'b0011100101100110;
    rom_data[3763]=16'b0111011001110000;
    rom_data[3764]=16'b0011100101010001;
    rom_data[3765]=16'b0111010101000100;
    rom_data[3766]=16'b0011100100111100;
    rom_data[3767]=16'b0111010000010110;
    rom_data[3768]=16'b0011100100100111;
    rom_data[3769]=16'b0111001011100101;
    rom_data[3770]=16'b0011100100010010;
    rom_data[3771]=16'b0111000110110001;
    rom_data[3772]=16'b0011100011111101;
    rom_data[3773]=16'b0111000001111100;
    rom_data[3774]=16'b0011100011101000;
    rom_data[3775]=16'b0110111101000100;
    rom_data[3776]=16'b0011100011010011;
    rom_data[3777]=16'b0110111000001011;
    rom_data[3778]=16'b0011100010111110;
    rom_data[3779]=16'b0110110011010000;
    rom_data[3780]=16'b0011100010101001;
    rom_data[3781]=16'b0110101110010011;
    rom_data[3782]=16'b0011100010010101;
    rom_data[3783]=16'b0110101001010101;
    rom_data[3784]=16'b0011100010000000;
    rom_data[3785]=16'b0110100100010110;
    rom_data[3786]=16'b0011100001101011;
    rom_data[3787]=16'b0110011111010101;
    rom_data[3788]=16'b0011100001010111;
    rom_data[3789]=16'b0110011010010100;
    rom_data[3790]=16'b0011100001000010;
    rom_data[3791]=16'b0110010101010010;
    rom_data[3792]=16'b0011100000101101;
    rom_data[3793]=16'b0110010000010000;
    rom_data[3794]=16'b0011100000011001;
    rom_data[3795]=16'b0110001011001100;
    rom_data[3796]=16'b0011100000000100;
    rom_data[3797]=16'b0110000110001001;
    rom_data[3798]=16'b0011011111101111;
    rom_data[3799]=16'b0110000001000101;
    rom_data[3800]=16'b0011011111011011;
    rom_data[3801]=16'b0101111100000001;
    rom_data[3802]=16'b0011011111000110;
    rom_data[3803]=16'b0101110110111100;
    rom_data[3804]=16'b0011011110110001;
    rom_data[3805]=16'b0101110001111000;
    rom_data[3806]=16'b0011011110011100;
    rom_data[3807]=16'b0101101100110100;
    rom_data[3808]=16'b0011011110000111;
    rom_data[3809]=16'b0101100111110001;
    rom_data[3810]=16'b0011011101110010;
    rom_data[3811]=16'b0101100010101110;
    rom_data[3812]=16'b0011011101011101;
    rom_data[3813]=16'b0101011101101011;
    rom_data[3814]=16'b0011011101001000;
    rom_data[3815]=16'b0101011000101001;
    rom_data[3816]=16'b0011011100110010;
    rom_data[3817]=16'b0101010011101000;
    rom_data[3818]=16'b0011011100011101;
    rom_data[3819]=16'b0101001110100111;
    rom_data[3820]=16'b0011011100000111;
    rom_data[3821]=16'b0101001001101000;
    rom_data[3822]=16'b0011011011110010;
    rom_data[3823]=16'b0101000100101010;
    rom_data[3824]=16'b0011011011011100;
    rom_data[3825]=16'b0100111111101101;
    rom_data[3826]=16'b0011011011000110;
    rom_data[3827]=16'b0100111010110010;
    rom_data[3828]=16'b0011011010110000;
    rom_data[3829]=16'b0100110101111000;
    rom_data[3830]=16'b0011011010011010;
    rom_data[3831]=16'b0100110001000000;
    rom_data[3832]=16'b0011011010000011;
    rom_data[3833]=16'b0100101100001010;
    rom_data[3834]=16'b0011011001101101;
    rom_data[3835]=16'b0100100111010110;
    rom_data[3836]=16'b0011011001010110;
    rom_data[3837]=16'b0100100010100101;
    rom_data[3838]=16'b0011011000111111;
    rom_data[3839]=16'b0100011101110110;
    rom_data[3840]=16'b0011011000101000;
    rom_data[3841]=16'b0100011001001001;
    rom_data[3842]=16'b0011011000010000;
    rom_data[3843]=16'b0100010100100000;
    rom_data[3844]=16'b0011010111111000;
    rom_data[3845]=16'b0100001111111001;
    rom_data[3846]=16'b0011010111100001;
    rom_data[3847]=16'b0100001011010110;
    rom_data[3848]=16'b0011010111001000;
    rom_data[3849]=16'b0100000110110111;
    rom_data[3850]=16'b0011010110110000;
    rom_data[3851]=16'b0100000010011100;
    rom_data[3852]=16'b0011010110010111;
    rom_data[3853]=16'b0011111110000100;
    rom_data[3854]=16'b0011010101111110;
    rom_data[3855]=16'b0011111001110010;
    rom_data[3856]=16'b0011010101100101;
    rom_data[3857]=16'b0011110101100100;
    rom_data[3858]=16'b0011010101001011;
    rom_data[3859]=16'b0011110001011011;
    rom_data[3860]=16'b0011010100110001;
    rom_data[3861]=16'b0011101101011000;
    rom_data[3862]=16'b0011010100010111;
    rom_data[3863]=16'b0011101001011011;
    rom_data[3864]=16'b0011010011111100;
    rom_data[3865]=16'b0011100101100100;
    rom_data[3866]=16'b0011010011100001;
    rom_data[3867]=16'b0011100001110100;
    rom_data[3868]=16'b0011010011000110;
    rom_data[3869]=16'b0011011110001100;
    rom_data[3870]=16'b0011010010101011;
    rom_data[3871]=16'b0011011010101100;
    rom_data[3872]=16'b0011010010001111;
    rom_data[3873]=16'b0011010111010100;
    rom_data[3874]=16'b0011010001110011;
    rom_data[3875]=16'b0011010100000101;
    rom_data[3876]=16'b0011010001010111;
    rom_data[3877]=16'b0011010000111111;
    rom_data[3878]=16'b0011010000111010;
    rom_data[3879]=16'b0011001110000101;
    rom_data[3880]=16'b0011010000011101;
    rom_data[3881]=16'b0011001011010101;
    rom_data[3882]=16'b0011010000000001;
    rom_data[3883]=16'b0011001000110001;
    rom_data[3884]=16'b0011001111100100;
    rom_data[3885]=16'b0011000110011001;
    rom_data[3886]=16'b0011001111000110;
    rom_data[3887]=16'b0011000100001111;
    rom_data[3888]=16'b0011001110101001;
    rom_data[3889]=16'b0011000010010010;
    rom_data[3890]=16'b0011001110001100;
    rom_data[3891]=16'b0011000000100100;
    rom_data[3892]=16'b0011001101101111;
    rom_data[3893]=16'b0010111111000101;
    rom_data[3894]=16'b0011001101010010;
    rom_data[3895]=16'b0010111101110110;
    rom_data[3896]=16'b0011001100110101;
    rom_data[3897]=16'b0010111100110111;
    rom_data[3898]=16'b0011001100011000;
    rom_data[3899]=16'b0010111100001001;
    rom_data[3900]=16'b0011001011111011;
    rom_data[3901]=16'b0010111011101100;
    rom_data[3902]=16'b0011001011011111;
    rom_data[3903]=16'b0010111011100000;
    rom_data[3904]=16'b0011001011000010;
    rom_data[3905]=16'b0010111011100110;
    rom_data[3906]=16'b0011001010100111;
    rom_data[3907]=16'b0010111011111110;
    rom_data[3908]=16'b0011001010001011;
    rom_data[3909]=16'b0010111100100110;
    rom_data[3910]=16'b0011001001101111;
    rom_data[3911]=16'b0010111101100000;
    rom_data[3912]=16'b0011001001010100;
    rom_data[3913]=16'b0010111110101011;
    rom_data[3914]=16'b0011001000111010;
    rom_data[3915]=16'b0011000000000110;
    rom_data[3916]=16'b0011001000011111;
    rom_data[3917]=16'b0011000001110000;
    rom_data[3918]=16'b0011001000000101;
    rom_data[3919]=16'b0011000011101010;
    rom_data[3920]=16'b0011000111101011;
    rom_data[3921]=16'b0011000101110010;
    rom_data[3922]=16'b0011000111010001;
    rom_data[3923]=16'b0011001000001000;
    rom_data[3924]=16'b0011000110111000;
    rom_data[3925]=16'b0011001010101010;
    rom_data[3926]=16'b0011000110011111;
    rom_data[3927]=16'b0011001101011001;
    rom_data[3928]=16'b0011000110000111;
    rom_data[3929]=16'b0011010000010100;
    rom_data[3930]=16'b0011000101101110;
    rom_data[3931]=16'b0011010011011001;
    rom_data[3932]=16'b0011000101010110;
    rom_data[3933]=16'b0011010110101000;
    rom_data[3934]=16'b0011000100111110;
    rom_data[3935]=16'b0011011010000001;
    rom_data[3936]=16'b0011000100100110;
    rom_data[3937]=16'b0011011101100011;
    rom_data[3938]=16'b0011000100001111;
    rom_data[3939]=16'b0011100001001100;
    rom_data[3940]=16'b0011000011111000;
    rom_data[3941]=16'b0011100100111110;
    rom_data[3942]=16'b0011000011100001;
    rom_data[3943]=16'b0011101000110110;
    rom_data[3944]=16'b0011000011001010;
    rom_data[3945]=16'b0011101100110101;
    rom_data[3946]=16'b0011000010110011;
    rom_data[3947]=16'b0011110000111010;
    rom_data[3948]=16'b0011000010011101;
    rom_data[3949]=16'b0011110101000101;
    rom_data[3950]=16'b0011000010000111;
    rom_data[3951]=16'b0011111001010101;
    rom_data[3952]=16'b0011000001110001;
    rom_data[3953]=16'b0011111101101010;
    rom_data[3954]=16'b0011000001011011;
    rom_data[3955]=16'b0100000010000011;
    rom_data[3956]=16'b0011000001000101;
    rom_data[3957]=16'b0100000110100001;
    rom_data[3958]=16'b0011000000101111;
    rom_data[3959]=16'b0100001011000011;
    rom_data[3960]=16'b0011000000011010;
    rom_data[3961]=16'b0100001111101000;
    rom_data[3962]=16'b0011000000000100;
    rom_data[3963]=16'b0100010100010000;
    rom_data[3964]=16'b0010111111101111;
    rom_data[3965]=16'b0100011000111100;
    rom_data[3966]=16'b0010111111011010;
    rom_data[3967]=16'b0100011101101010;
    rom_data[3968]=16'b0010111111000101;
    rom_data[3969]=16'b0100100010011011;
    rom_data[3970]=16'b0010111110110000;
    rom_data[3971]=16'b0100100111001111;
    rom_data[3972]=16'b0010111110011011;
    rom_data[3973]=16'b0100101100000100;
    rom_data[3974]=16'b0010111110000110;
    rom_data[3975]=16'b0100110000111100;
    rom_data[3976]=16'b0010111101110001;
    rom_data[3977]=16'b0100110101110101;
    rom_data[3978]=16'b0010111101011100;
    rom_data[3979]=16'b0100111010110001;
    rom_data[3980]=16'b0010111101000111;
    rom_data[3981]=16'b0100111111101101;
    rom_data[3982]=16'b0010111100110011;
    rom_data[3983]=16'b0101000100101011;
    rom_data[3984]=16'b0010111100011110;
    rom_data[3985]=16'b0101001001101010;
    rom_data[3986]=16'b0010111100001001;
    rom_data[3987]=16'b0101001110101011;
    rom_data[3988]=16'b0010111011110101;
    rom_data[3989]=16'b0101010011101100;
    rom_data[3990]=16'b0010111011100000;
    rom_data[3991]=16'b0101011000101110;
    rom_data[3992]=16'b0010111011100000;
    rom_data[3993]=16'b0101011101110001;
    rom_data[3994]=16'b0010111011110101;
    rom_data[3995]=16'b0101100010110100;
    rom_data[3996]=16'b0010111100001001;
    rom_data[3997]=16'b0101100111110111;
    rom_data[3998]=16'b0010111100011110;
    rom_data[3999]=16'b0101101100111011;
    rom_data[4000]=16'b0010111100110011;
    rom_data[4001]=16'b0101110010000000;





    if (addr[0]==1'b0) begin
        data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
    end else begin //data in 50%
        
        case (addr[2:1])
            2'b00: begin // this is a CHANNEL A
                data_d = {6'b000110, addr[2:1], CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                data_d = {6'b000110, addr[2:1], CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                data_d = {6'b000110, addr[2:1], CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                data_d = {6'b000110, addr[2:1], CH_D_q};
            end

            default: begin
            end
        endcase

    end // if VREF
end // always


always @(posedge addr[0]) begin
    CH_A_q<=CH_A_d;
    CH_B_q<=CH_B_d;
    CH_C_q<=CH_C_d;
    CH_D_q<=CH_D_d;
end


always @(posedge clk) begin
  if (addr==0) begin
    data_q <= 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (addr==1) begin
    data_q <= 24'b00111000_0000000000000000;    // set Vref only once
  end else begin
    data_q <= data_d;
  end
end // always
 
endmodule