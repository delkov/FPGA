module mems_rom_9 (
    input clk,
    input [8:0] addr,
    // input [7:0] delta_A,
    // input [7:0] delta_B,
    // input [7:0] delta_C,
    // input [7:0] delta_D,
    output [23:0] data
  );
 
  reg [23:0] rom_data [481:0];
  reg [23:0] data_d, data_q;
 
  assign data = data_q;
 
  always @(*) begin

  // OLDVI STYLE
  // rom_data[0] = 24'b001010000000000000000001; // SOFT_RESET;
  // rom_data[1] = 24'b001101110011111111111111;//1111; // LDAC SETUP

  // rom_data[2] = {8'b00010000, delta_A, 8'b00011111}; // CH A
  // rom_data[3] = {8'b00010001, delta_B, 8'b00000000}; // CH B
  // rom_data[4] = {8'b00010010, delta_C, 8'b00011111}; // CH C
  // rom_data[5] = {8'b00010011, delta_D, 8'b00000000}; // CH D

  // NEW
    rom_data[0] = 24'b001010000000000000000001; // SOFT_RESET;
    rom_data[1] = 24'b001101110011111111110000;//1111; // LDAC SETUP

    // rom_data[2] = {8'b00000000, delta_A, 8'b00000000}; // CH A
    // rom_data[3] = {8'b00000001, delta_B, 8'b00000000}; // CH B
    // rom_data[4] = {8'b00000010, delta_C, 8'b00000000}; // CH C
    // rom_data[5] = {8'b00010011, delta_D, 8'b00000000}; // CH D

    rom_data[2]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[6]={8'b00000000,8'b01011101,8'b00000000};
    rom_data[10]={8'b00000000,8'b01101001,8'b00000000};
    rom_data[14]={8'b00000000,8'b01110100,8'b00000000};
    rom_data[18]={8'b00000000,8'b01111110,8'b00000000};
    rom_data[22]={8'b00000000,8'b10000101,8'b00000000};
    rom_data[26]={8'b00000000,8'b10001010,8'b00000000};
    rom_data[30]={8'b00000000,8'b10001100,8'b00000000};
    rom_data[34]={8'b00000000,8'b10001011,8'b00000000};
    rom_data[38]={8'b00000000,8'b10001000,8'b00000000};
    rom_data[42]={8'b00000000,8'b10000010,8'b00000000};
    rom_data[46]={8'b00000000,8'b01111001,8'b00000000};
    rom_data[50]={8'b00000000,8'b01101111,8'b00000000};
    rom_data[54]={8'b00000000,8'b01100011,8'b00000000};
    rom_data[58]={8'b00000000,8'b01010110,8'b00000000};
    rom_data[62]={8'b00000000,8'b01001010,8'b00000000};
    rom_data[66]={8'b00000000,8'b00111101,8'b00000000};
    rom_data[70]={8'b00000000,8'b00110001,8'b00000000};
    rom_data[74]={8'b00000000,8'b00100111,8'b00000000};
    rom_data[78]={8'b00000000,8'b00011110,8'b00000000};
    rom_data[82]={8'b00000000,8'b00011000,8'b00000000};
    rom_data[86]={8'b00000000,8'b00010101,8'b00000000};
    rom_data[90]={8'b00000000,8'b00010100,8'b00000000};
    rom_data[94]={8'b00000000,8'b00010110,8'b00000000};
    rom_data[98]={8'b00000000,8'b00011011,8'b00000000};
    rom_data[102]={8'b00000000,8'b00100010,8'b00000000};
    rom_data[106]={8'b00000000,8'b00101100,8'b00000000};
    rom_data[110]={8'b00000000,8'b00110111,8'b00000000};
    rom_data[114]={8'b00000000,8'b01000011,8'b00000000};
    rom_data[118]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[122]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[126]={8'b00000000,8'b01011101,8'b00000000};
    rom_data[130]={8'b00000000,8'b01101001,8'b00000000};
    rom_data[134]={8'b00000000,8'b01110100,8'b00000000};
    rom_data[138]={8'b00000000,8'b01111110,8'b00000000};
    rom_data[142]={8'b00000000,8'b10000101,8'b00000000};
    rom_data[146]={8'b00000000,8'b10001010,8'b00000000};
    rom_data[150]={8'b00000000,8'b10001100,8'b00000000};
    rom_data[154]={8'b00000000,8'b10001011,8'b00000000};
    rom_data[158]={8'b00000000,8'b10001000,8'b00000000};
    rom_data[162]={8'b00000000,8'b10000010,8'b00000000};
    rom_data[166]={8'b00000000,8'b01111001,8'b00000000};
    rom_data[170]={8'b00000000,8'b01101111,8'b00000000};
    rom_data[174]={8'b00000000,8'b01100011,8'b00000000};
    rom_data[178]={8'b00000000,8'b01010110,8'b00000000};
    rom_data[182]={8'b00000000,8'b01001010,8'b00000000};
    rom_data[186]={8'b00000000,8'b00111101,8'b00000000};
    rom_data[190]={8'b00000000,8'b00110001,8'b00000000};
    rom_data[194]={8'b00000000,8'b00100111,8'b00000000};
    rom_data[198]={8'b00000000,8'b00011110,8'b00000000};
    rom_data[202]={8'b00000000,8'b00011000,8'b00000000};
    rom_data[206]={8'b00000000,8'b00010101,8'b00000000};
    rom_data[210]={8'b00000000,8'b00010100,8'b00000000};
    rom_data[214]={8'b00000000,8'b00010110,8'b00000000};
    rom_data[218]={8'b00000000,8'b00011011,8'b00000000};
    rom_data[222]={8'b00000000,8'b00100010,8'b00000000};
    rom_data[226]={8'b00000000,8'b00101100,8'b00000000};
    rom_data[230]={8'b00000000,8'b00110111,8'b00000000};
    rom_data[234]={8'b00000000,8'b01000011,8'b00000000};
    rom_data[238]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[242]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[246]={8'b00000000,8'b01011101,8'b00000000};
    rom_data[250]={8'b00000000,8'b01101001,8'b00000000};
    rom_data[254]={8'b00000000,8'b01110100,8'b00000000};
    rom_data[258]={8'b00000000,8'b01111110,8'b00000000};
    rom_data[262]={8'b00000000,8'b10000101,8'b00000000};
    rom_data[266]={8'b00000000,8'b10001010,8'b00000000};
    rom_data[270]={8'b00000000,8'b10001100,8'b00000000};
    rom_data[274]={8'b00000000,8'b10001011,8'b00000000};
    rom_data[278]={8'b00000000,8'b10001000,8'b00000000};
    rom_data[282]={8'b00000000,8'b10000010,8'b00000000};
    rom_data[286]={8'b00000000,8'b01111001,8'b00000000};
    rom_data[290]={8'b00000000,8'b01101111,8'b00000000};
    rom_data[294]={8'b00000000,8'b01100011,8'b00000000};
    rom_data[298]={8'b00000000,8'b01010110,8'b00000000};
    rom_data[302]={8'b00000000,8'b01001010,8'b00000000};
    rom_data[306]={8'b00000000,8'b00111101,8'b00000000};
    rom_data[310]={8'b00000000,8'b00110001,8'b00000000};
    rom_data[314]={8'b00000000,8'b00100111,8'b00000000};
    rom_data[318]={8'b00000000,8'b00011110,8'b00000000};
    rom_data[322]={8'b00000000,8'b00011000,8'b00000000};
    rom_data[326]={8'b00000000,8'b00010101,8'b00000000};
    rom_data[330]={8'b00000000,8'b00010100,8'b00000000};
    rom_data[334]={8'b00000000,8'b00010110,8'b00000000};
    rom_data[338]={8'b00000000,8'b00011011,8'b00000000};
    rom_data[342]={8'b00000000,8'b00100010,8'b00000000};
    rom_data[346]={8'b00000000,8'b00101100,8'b00000000};
    rom_data[350]={8'b00000000,8'b00110111,8'b00000000};
    rom_data[354]={8'b00000000,8'b01000011,8'b00000000};
    rom_data[358]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[362]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[366]={8'b00000000,8'b01011101,8'b00000000};
    rom_data[370]={8'b00000000,8'b01101001,8'b00000000};
    rom_data[374]={8'b00000000,8'b01110100,8'b00000000};
    rom_data[378]={8'b00000000,8'b01111110,8'b00000000};
    rom_data[382]={8'b00000000,8'b10000101,8'b00000000};
    rom_data[386]={8'b00000000,8'b10001010,8'b00000000};
    rom_data[390]={8'b00000000,8'b10001100,8'b00000000};
    rom_data[394]={8'b00000000,8'b10001011,8'b00000000};
    rom_data[398]={8'b00000000,8'b10001000,8'b00000000};
    rom_data[402]={8'b00000000,8'b10000010,8'b00000000};
    rom_data[406]={8'b00000000,8'b01111001,8'b00000000};
    rom_data[410]={8'b00000000,8'b01101111,8'b00000000};
    rom_data[414]={8'b00000000,8'b01100011,8'b00000000};
    rom_data[418]={8'b00000000,8'b01010110,8'b00000000};
    rom_data[422]={8'b00000000,8'b01001010,8'b00000000};
    rom_data[426]={8'b00000000,8'b00111101,8'b00000000};
    rom_data[430]={8'b00000000,8'b00110001,8'b00000000};
    rom_data[434]={8'b00000000,8'b00100111,8'b00000000};
    rom_data[438]={8'b00000000,8'b00011110,8'b00000000};
    rom_data[442]={8'b00000000,8'b00011000,8'b00000000};
    rom_data[446]={8'b00000000,8'b00010101,8'b00000000};
    rom_data[450]={8'b00000000,8'b00010100,8'b00000000};
    rom_data[454]={8'b00000000,8'b00010110,8'b00000000};
    rom_data[458]={8'b00000000,8'b00011011,8'b00000000};
    rom_data[462]={8'b00000000,8'b00100010,8'b00000000};
    rom_data[466]={8'b00000000,8'b00101100,8'b00000000};
    rom_data[470]={8'b00000000,8'b00110111,8'b00000000};
    rom_data[474]={8'b00000000,8'b01000011,8'b00000000};
    rom_data[478]={8'b00000000,8'b01010000,8'b00000000};
    rom_data[3]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[7]={8'b00000001,8'b01000011,8'b00000000};
    rom_data[11]={8'b00000001,8'b00110111,8'b00000000};
    rom_data[15]={8'b00000001,8'b00101100,8'b00000000};
    rom_data[19]={8'b00000001,8'b00100010,8'b00000000};
    rom_data[23]={8'b00000001,8'b00011011,8'b00000000};
    rom_data[27]={8'b00000001,8'b00010110,8'b00000000};
    rom_data[31]={8'b00000001,8'b00010100,8'b00000000};
    rom_data[35]={8'b00000001,8'b00010101,8'b00000000};
    rom_data[39]={8'b00000001,8'b00011000,8'b00000000};
    rom_data[43]={8'b00000001,8'b00011110,8'b00000000};
    rom_data[47]={8'b00000001,8'b00100111,8'b00000000};
    rom_data[51]={8'b00000001,8'b00110001,8'b00000000};
    rom_data[55]={8'b00000001,8'b00111101,8'b00000000};
    rom_data[59]={8'b00000001,8'b01001010,8'b00000000};
    rom_data[63]={8'b00000001,8'b01010110,8'b00000000};
    rom_data[67]={8'b00000001,8'b01100011,8'b00000000};
    rom_data[71]={8'b00000001,8'b01101111,8'b00000000};
    rom_data[75]={8'b00000001,8'b01111001,8'b00000000};
    rom_data[79]={8'b00000001,8'b10000010,8'b00000000};
    rom_data[83]={8'b00000001,8'b10001000,8'b00000000};
    rom_data[87]={8'b00000001,8'b10001011,8'b00000000};
    rom_data[91]={8'b00000001,8'b10001100,8'b00000000};
    rom_data[95]={8'b00000001,8'b10001010,8'b00000000};
    rom_data[99]={8'b00000001,8'b10000101,8'b00000000};
    rom_data[103]={8'b00000001,8'b01111110,8'b00000000};
    rom_data[107]={8'b00000001,8'b01110100,8'b00000000};
    rom_data[111]={8'b00000001,8'b01101001,8'b00000000};
    rom_data[115]={8'b00000001,8'b01011101,8'b00000000};
    rom_data[119]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[123]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[127]={8'b00000001,8'b01000011,8'b00000000};
    rom_data[131]={8'b00000001,8'b00110111,8'b00000000};
    rom_data[135]={8'b00000001,8'b00101100,8'b00000000};
    rom_data[139]={8'b00000001,8'b00100010,8'b00000000};
    rom_data[143]={8'b00000001,8'b00011011,8'b00000000};
    rom_data[147]={8'b00000001,8'b00010110,8'b00000000};
    rom_data[151]={8'b00000001,8'b00010100,8'b00000000};
    rom_data[155]={8'b00000001,8'b00010101,8'b00000000};
    rom_data[159]={8'b00000001,8'b00011000,8'b00000000};
    rom_data[163]={8'b00000001,8'b00011110,8'b00000000};
    rom_data[167]={8'b00000001,8'b00100111,8'b00000000};
    rom_data[171]={8'b00000001,8'b00110001,8'b00000000};
    rom_data[175]={8'b00000001,8'b00111101,8'b00000000};
    rom_data[179]={8'b00000001,8'b01001010,8'b00000000};
    rom_data[183]={8'b00000001,8'b01010110,8'b00000000};
    rom_data[187]={8'b00000001,8'b01100011,8'b00000000};
    rom_data[191]={8'b00000001,8'b01101111,8'b00000000};
    rom_data[195]={8'b00000001,8'b01111001,8'b00000000};
    rom_data[199]={8'b00000001,8'b10000010,8'b00000000};
    rom_data[203]={8'b00000001,8'b10001000,8'b00000000};
    rom_data[207]={8'b00000001,8'b10001011,8'b00000000};
    rom_data[211]={8'b00000001,8'b10001100,8'b00000000};
    rom_data[215]={8'b00000001,8'b10001010,8'b00000000};
    rom_data[219]={8'b00000001,8'b10000101,8'b00000000};
    rom_data[223]={8'b00000001,8'b01111110,8'b00000000};
    rom_data[227]={8'b00000001,8'b01110100,8'b00000000};
    rom_data[231]={8'b00000001,8'b01101001,8'b00000000};
    rom_data[235]={8'b00000001,8'b01011101,8'b00000000};
    rom_data[239]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[243]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[247]={8'b00000001,8'b01000011,8'b00000000};
    rom_data[251]={8'b00000001,8'b00110111,8'b00000000};
    rom_data[255]={8'b00000001,8'b00101100,8'b00000000};
    rom_data[259]={8'b00000001,8'b00100010,8'b00000000};
    rom_data[263]={8'b00000001,8'b00011011,8'b00000000};
    rom_data[267]={8'b00000001,8'b00010110,8'b00000000};
    rom_data[271]={8'b00000001,8'b00010100,8'b00000000};
    rom_data[275]={8'b00000001,8'b00010101,8'b00000000};
    rom_data[279]={8'b00000001,8'b00011000,8'b00000000};
    rom_data[283]={8'b00000001,8'b00011110,8'b00000000};
    rom_data[287]={8'b00000001,8'b00100111,8'b00000000};
    rom_data[291]={8'b00000001,8'b00110001,8'b00000000};
    rom_data[295]={8'b00000001,8'b00111101,8'b00000000};
    rom_data[299]={8'b00000001,8'b01001010,8'b00000000};
    rom_data[303]={8'b00000001,8'b01010110,8'b00000000};
    rom_data[307]={8'b00000001,8'b01100011,8'b00000000};
    rom_data[311]={8'b00000001,8'b01101111,8'b00000000};
    rom_data[315]={8'b00000001,8'b01111001,8'b00000000};
    rom_data[319]={8'b00000001,8'b10000010,8'b00000000};
    rom_data[323]={8'b00000001,8'b10001000,8'b00000000};
    rom_data[327]={8'b00000001,8'b10001011,8'b00000000};
    rom_data[331]={8'b00000001,8'b10001100,8'b00000000};
    rom_data[335]={8'b00000001,8'b10001010,8'b00000000};
    rom_data[339]={8'b00000001,8'b10000101,8'b00000000};
    rom_data[343]={8'b00000001,8'b01111110,8'b00000000};
    rom_data[347]={8'b00000001,8'b01110100,8'b00000000};
    rom_data[351]={8'b00000001,8'b01101001,8'b00000000};
    rom_data[355]={8'b00000001,8'b01011101,8'b00000000};
    rom_data[359]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[363]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[367]={8'b00000001,8'b01000011,8'b00000000};
    rom_data[371]={8'b00000001,8'b00110111,8'b00000000};
    rom_data[375]={8'b00000001,8'b00101100,8'b00000000};
    rom_data[379]={8'b00000001,8'b00100010,8'b00000000};
    rom_data[383]={8'b00000001,8'b00011011,8'b00000000};
    rom_data[387]={8'b00000001,8'b00010110,8'b00000000};
    rom_data[391]={8'b00000001,8'b00010100,8'b00000000};
    rom_data[395]={8'b00000001,8'b00010101,8'b00000000};
    rom_data[399]={8'b00000001,8'b00011000,8'b00000000};
    rom_data[403]={8'b00000001,8'b00011110,8'b00000000};
    rom_data[407]={8'b00000001,8'b00100111,8'b00000000};
    rom_data[411]={8'b00000001,8'b00110001,8'b00000000};
    rom_data[415]={8'b00000001,8'b00111101,8'b00000000};
    rom_data[419]={8'b00000001,8'b01001010,8'b00000000};
    rom_data[423]={8'b00000001,8'b01010110,8'b00000000};
    rom_data[427]={8'b00000001,8'b01100011,8'b00000000};
    rom_data[431]={8'b00000001,8'b01101111,8'b00000000};
    rom_data[435]={8'b00000001,8'b01111001,8'b00000000};
    rom_data[439]={8'b00000001,8'b10000010,8'b00000000};
    rom_data[443]={8'b00000001,8'b10001000,8'b00000000};
    rom_data[447]={8'b00000001,8'b10001011,8'b00000000};
    rom_data[451]={8'b00000001,8'b10001100,8'b00000000};
    rom_data[455]={8'b00000001,8'b10001010,8'b00000000};
    rom_data[459]={8'b00000001,8'b10000101,8'b00000000};
    rom_data[463]={8'b00000001,8'b01111110,8'b00000000};
    rom_data[467]={8'b00000001,8'b01110100,8'b00000000};
    rom_data[471]={8'b00000001,8'b01101001,8'b00000000};
    rom_data[475]={8'b00000001,8'b01011101,8'b00000000};
    rom_data[479]={8'b00000001,8'b01010000,8'b00000000};
    rom_data[4]={8'b00000010,8'b00010100,8'b00000000};
    rom_data[8]={8'b00000010,8'b00010101,8'b00000000};
    rom_data[12]={8'b00000010,8'b00010110,8'b00000000};
    rom_data[16]={8'b00000010,8'b00010111,8'b00000000};
    rom_data[20]={8'b00000010,8'b00011000,8'b00000000};
    rom_data[24]={8'b00000010,8'b00011001,8'b00000000};
    rom_data[28]={8'b00000010,8'b00011010,8'b00000000};
    rom_data[32]={8'b00000010,8'b00011011,8'b00000000};
    rom_data[36]={8'b00000010,8'b00011100,8'b00000000};
    rom_data[40]={8'b00000010,8'b00011101,8'b00000000};
    rom_data[44]={8'b00000010,8'b00011110,8'b00000000};
    rom_data[48]={8'b00000010,8'b00011111,8'b00000000};
    rom_data[52]={8'b00000010,8'b00100000,8'b00000000};
    rom_data[56]={8'b00000010,8'b00100001,8'b00000000};
    rom_data[60]={8'b00000010,8'b00100010,8'b00000000};
    rom_data[64]={8'b00000010,8'b00100011,8'b00000000};
    rom_data[68]={8'b00000010,8'b00100100,8'b00000000};
    rom_data[72]={8'b00000010,8'b00100101,8'b00000000};
    rom_data[76]={8'b00000010,8'b00100110,8'b00000000};
    rom_data[80]={8'b00000010,8'b00100111,8'b00000000};
    rom_data[84]={8'b00000010,8'b00101000,8'b00000000};
    rom_data[88]={8'b00000010,8'b00101001,8'b00000000};
    rom_data[92]={8'b00000010,8'b00101010,8'b00000000};
    rom_data[96]={8'b00000010,8'b00101011,8'b00000000};
    rom_data[100]={8'b00000010,8'b00101100,8'b00000000};
    rom_data[104]={8'b00000010,8'b00101101,8'b00000000};
    rom_data[108]={8'b00000010,8'b00101110,8'b00000000};
    rom_data[112]={8'b00000010,8'b00101111,8'b00000000};
    rom_data[116]={8'b00000010,8'b00110000,8'b00000000};
    rom_data[120]={8'b00000010,8'b00110001,8'b00000000};
    rom_data[124]={8'b00000010,8'b00110010,8'b00000000};
    rom_data[128]={8'b00000010,8'b00110011,8'b00000000};
    rom_data[132]={8'b00000010,8'b00110100,8'b00000000};
    rom_data[136]={8'b00000010,8'b00110101,8'b00000000};
    rom_data[140]={8'b00000010,8'b00110110,8'b00000000};
    rom_data[144]={8'b00000010,8'b00110111,8'b00000000};
    rom_data[148]={8'b00000010,8'b00111000,8'b00000000};
    rom_data[152]={8'b00000010,8'b00111001,8'b00000000};
    rom_data[156]={8'b00000010,8'b00111010,8'b00000000};
    rom_data[160]={8'b00000010,8'b00111011,8'b00000000};
    rom_data[164]={8'b00000010,8'b00111100,8'b00000000};
    rom_data[168]={8'b00000010,8'b00111101,8'b00000000};
    rom_data[172]={8'b00000010,8'b00111110,8'b00000000};
    rom_data[176]={8'b00000010,8'b00111111,8'b00000000};
    rom_data[180]={8'b00000010,8'b01000000,8'b00000000};
    rom_data[184]={8'b00000010,8'b01000001,8'b00000000};
    rom_data[188]={8'b00000010,8'b01000010,8'b00000000};
    rom_data[192]={8'b00000010,8'b01000011,8'b00000000};
    rom_data[196]={8'b00000010,8'b01000100,8'b00000000};
    rom_data[200]={8'b00000010,8'b01000101,8'b00000000};
    rom_data[204]={8'b00000010,8'b01000110,8'b00000000};
    rom_data[208]={8'b00000010,8'b01000111,8'b00000000};
    rom_data[212]={8'b00000010,8'b01001000,8'b00000000};
    rom_data[216]={8'b00000010,8'b01001001,8'b00000000};
    rom_data[220]={8'b00000010,8'b01001010,8'b00000000};
    rom_data[224]={8'b00000010,8'b01001011,8'b00000000};
    rom_data[228]={8'b00000010,8'b01001100,8'b00000000};
    rom_data[232]={8'b00000010,8'b01001101,8'b00000000};
    rom_data[236]={8'b00000010,8'b01001110,8'b00000000};
    rom_data[240]={8'b00000010,8'b01001111,8'b00000000};
    rom_data[244]={8'b00000010,8'b01010001,8'b00000000};
    rom_data[248]={8'b00000010,8'b01010010,8'b00000000};
    rom_data[252]={8'b00000010,8'b01010011,8'b00000000};
    rom_data[256]={8'b00000010,8'b01010100,8'b00000000};
    rom_data[260]={8'b00000010,8'b01010101,8'b00000000};
    rom_data[264]={8'b00000010,8'b01010110,8'b00000000};
    rom_data[268]={8'b00000010,8'b01010111,8'b00000000};
    rom_data[272]={8'b00000010,8'b01011000,8'b00000000};
    rom_data[276]={8'b00000010,8'b01011001,8'b00000000};
    rom_data[280]={8'b00000010,8'b01011010,8'b00000000};
    rom_data[284]={8'b00000010,8'b01011011,8'b00000000};
    rom_data[288]={8'b00000010,8'b01011100,8'b00000000};
    rom_data[292]={8'b00000010,8'b01011101,8'b00000000};
    rom_data[296]={8'b00000010,8'b01011110,8'b00000000};
    rom_data[300]={8'b00000010,8'b01011111,8'b00000000};
    rom_data[304]={8'b00000010,8'b01100000,8'b00000000};
    rom_data[308]={8'b00000010,8'b01100001,8'b00000000};
    rom_data[312]={8'b00000010,8'b01100010,8'b00000000};
    rom_data[316]={8'b00000010,8'b01100011,8'b00000000};
    rom_data[320]={8'b00000010,8'b01100100,8'b00000000};
    rom_data[324]={8'b00000010,8'b01100101,8'b00000000};
    rom_data[328]={8'b00000010,8'b01100110,8'b00000000};
    rom_data[332]={8'b00000010,8'b01100111,8'b00000000};
    rom_data[336]={8'b00000010,8'b01101000,8'b00000000};
    rom_data[340]={8'b00000010,8'b01101001,8'b00000000};
    rom_data[344]={8'b00000010,8'b01101010,8'b00000000};
    rom_data[348]={8'b00000010,8'b01101011,8'b00000000};
    rom_data[352]={8'b00000010,8'b01101100,8'b00000000};
    rom_data[356]={8'b00000010,8'b01101101,8'b00000000};
    rom_data[360]={8'b00000010,8'b01101110,8'b00000000};
    rom_data[364]={8'b00000010,8'b01101111,8'b00000000};
    rom_data[368]={8'b00000010,8'b01110000,8'b00000000};
    rom_data[372]={8'b00000010,8'b01110001,8'b00000000};
    rom_data[376]={8'b00000010,8'b01110010,8'b00000000};
    rom_data[380]={8'b00000010,8'b01110011,8'b00000000};
    rom_data[384]={8'b00000010,8'b01110100,8'b00000000};
    rom_data[388]={8'b00000010,8'b01110101,8'b00000000};
    rom_data[392]={8'b00000010,8'b01110110,8'b00000000};
    rom_data[396]={8'b00000010,8'b01110111,8'b00000000};
    rom_data[400]={8'b00000010,8'b01111000,8'b00000000};
    rom_data[404]={8'b00000010,8'b01111001,8'b00000000};
    rom_data[408]={8'b00000010,8'b01111010,8'b00000000};
    rom_data[412]={8'b00000010,8'b01111011,8'b00000000};
    rom_data[416]={8'b00000010,8'b01111100,8'b00000000};
    rom_data[420]={8'b00000010,8'b01111101,8'b00000000};
    rom_data[424]={8'b00000010,8'b01111110,8'b00000000};
    rom_data[428]={8'b00000010,8'b01111111,8'b00000000};
    rom_data[432]={8'b00000010,8'b10000000,8'b00000000};
    rom_data[436]={8'b00000010,8'b10000001,8'b00000000};
    rom_data[440]={8'b00000010,8'b10000010,8'b00000000};
    rom_data[444]={8'b00000010,8'b10000011,8'b00000000};
    rom_data[448]={8'b00000010,8'b10000100,8'b00000000};
    rom_data[452]={8'b00000010,8'b10000101,8'b00000000};
    rom_data[456]={8'b00000010,8'b10000110,8'b00000000};
    rom_data[460]={8'b00000010,8'b10000111,8'b00000000};
    rom_data[464]={8'b00000010,8'b10001000,8'b00000000};
    rom_data[468]={8'b00000010,8'b10001001,8'b00000000};
    rom_data[472]={8'b00000010,8'b10001010,8'b00000000};
    rom_data[476]={8'b00000010,8'b10001011,8'b00000000};
    rom_data[480]={8'b00000010,8'b10001100,8'b00000000};
    rom_data[5]={8'b00010011,8'b10001100,8'b00000000};
    rom_data[9]={8'b00010011,8'b10001011,8'b00000000};
    rom_data[13]={8'b00010011,8'b10001010,8'b00000000};
    rom_data[17]={8'b00010011,8'b10001001,8'b00000000};
    rom_data[21]={8'b00010011,8'b10001000,8'b00000000};
    rom_data[25]={8'b00010011,8'b10000111,8'b00000000};
    rom_data[29]={8'b00010011,8'b10000110,8'b00000000};
    rom_data[33]={8'b00010011,8'b10000101,8'b00000000};
    rom_data[37]={8'b00010011,8'b10000100,8'b00000000};
    rom_data[41]={8'b00010011,8'b10000011,8'b00000000};
    rom_data[45]={8'b00010011,8'b10000010,8'b00000000};
    rom_data[49]={8'b00010011,8'b10000001,8'b00000000};
    rom_data[53]={8'b00010011,8'b10000000,8'b00000000};
    rom_data[57]={8'b00010011,8'b01111111,8'b00000000};
    rom_data[61]={8'b00010011,8'b01111110,8'b00000000};
    rom_data[65]={8'b00010011,8'b01111101,8'b00000000};
    rom_data[69]={8'b00010011,8'b01111100,8'b00000000};
    rom_data[73]={8'b00010011,8'b01111011,8'b00000000};
    rom_data[77]={8'b00010011,8'b01111010,8'b00000000};
    rom_data[81]={8'b00010011,8'b01111001,8'b00000000};
    rom_data[85]={8'b00010011,8'b01111000,8'b00000000};
    rom_data[89]={8'b00010011,8'b01110111,8'b00000000};
    rom_data[93]={8'b00010011,8'b01110110,8'b00000000};
    rom_data[97]={8'b00010011,8'b01110101,8'b00000000};
    rom_data[101]={8'b00010011,8'b01110100,8'b00000000};
    rom_data[105]={8'b00010011,8'b01110011,8'b00000000};
    rom_data[109]={8'b00010011,8'b01110010,8'b00000000};
    rom_data[113]={8'b00010011,8'b01110001,8'b00000000};
    rom_data[117]={8'b00010011,8'b01110000,8'b00000000};
    rom_data[121]={8'b00010011,8'b01101111,8'b00000000};
    rom_data[125]={8'b00010011,8'b01101110,8'b00000000};
    rom_data[129]={8'b00010011,8'b01101101,8'b00000000};
    rom_data[133]={8'b00010011,8'b01101100,8'b00000000};
    rom_data[137]={8'b00010011,8'b01101011,8'b00000000};
    rom_data[141]={8'b00010011,8'b01101010,8'b00000000};
    rom_data[145]={8'b00010011,8'b01101001,8'b00000000};
    rom_data[149]={8'b00010011,8'b01101000,8'b00000000};
    rom_data[153]={8'b00010011,8'b01100111,8'b00000000};
    rom_data[157]={8'b00010011,8'b01100110,8'b00000000};
    rom_data[161]={8'b00010011,8'b01100101,8'b00000000};
    rom_data[165]={8'b00010011,8'b01100100,8'b00000000};
    rom_data[169]={8'b00010011,8'b01100011,8'b00000000};
    rom_data[173]={8'b00010011,8'b01100010,8'b00000000};
    rom_data[177]={8'b00010011,8'b01100001,8'b00000000};
    rom_data[181]={8'b00010011,8'b01100000,8'b00000000};
    rom_data[185]={8'b00010011,8'b01011111,8'b00000000};
    rom_data[189]={8'b00010011,8'b01011110,8'b00000000};
    rom_data[193]={8'b00010011,8'b01011101,8'b00000000};
    rom_data[197]={8'b00010011,8'b01011100,8'b00000000};
    rom_data[201]={8'b00010011,8'b01011011,8'b00000000};
    rom_data[205]={8'b00010011,8'b01011010,8'b00000000};
    rom_data[209]={8'b00010011,8'b01011001,8'b00000000};
    rom_data[213]={8'b00010011,8'b01011000,8'b00000000};
    rom_data[217]={8'b00010011,8'b01010111,8'b00000000};
    rom_data[221]={8'b00010011,8'b01010110,8'b00000000};
    rom_data[225]={8'b00010011,8'b01010101,8'b00000000};
    rom_data[229]={8'b00010011,8'b01010100,8'b00000000};
    rom_data[233]={8'b00010011,8'b01010011,8'b00000000};
    rom_data[237]={8'b00010011,8'b01010010,8'b00000000};
    rom_data[241]={8'b00010011,8'b01010001,8'b00000000};
    rom_data[245]={8'b00010011,8'b01001111,8'b00000000};
    rom_data[249]={8'b00010011,8'b01001110,8'b00000000};
    rom_data[253]={8'b00010011,8'b01001101,8'b00000000};
    rom_data[257]={8'b00010011,8'b01001100,8'b00000000};
    rom_data[261]={8'b00010011,8'b01001011,8'b00000000};
    rom_data[265]={8'b00010011,8'b01001010,8'b00000000};
    rom_data[269]={8'b00010011,8'b01001001,8'b00000000};
    rom_data[273]={8'b00010011,8'b01001000,8'b00000000};
    rom_data[277]={8'b00010011,8'b01000111,8'b00000000};
    rom_data[281]={8'b00010011,8'b01000110,8'b00000000};
    rom_data[285]={8'b00010011,8'b01000101,8'b00000000};
    rom_data[289]={8'b00010011,8'b01000100,8'b00000000};
    rom_data[293]={8'b00010011,8'b01000011,8'b00000000};
    rom_data[297]={8'b00010011,8'b01000010,8'b00000000};
    rom_data[301]={8'b00010011,8'b01000001,8'b00000000};
    rom_data[305]={8'b00010011,8'b01000000,8'b00000000};
    rom_data[309]={8'b00010011,8'b00111111,8'b00000000};
    rom_data[313]={8'b00010011,8'b00111110,8'b00000000};
    rom_data[317]={8'b00010011,8'b00111101,8'b00000000};
    rom_data[321]={8'b00010011,8'b00111100,8'b00000000};
    rom_data[325]={8'b00010011,8'b00111011,8'b00000000};
    rom_data[329]={8'b00010011,8'b00111010,8'b00000000};
    rom_data[333]={8'b00010011,8'b00111001,8'b00000000};
    rom_data[337]={8'b00010011,8'b00111000,8'b00000000};
    rom_data[341]={8'b00010011,8'b00110111,8'b00000000};
    rom_data[345]={8'b00010011,8'b00110110,8'b00000000};
    rom_data[349]={8'b00010011,8'b00110101,8'b00000000};
    rom_data[353]={8'b00010011,8'b00110100,8'b00000000};
    rom_data[357]={8'b00010011,8'b00110011,8'b00000000};
    rom_data[361]={8'b00010011,8'b00110010,8'b00000000};
    rom_data[365]={8'b00010011,8'b00110001,8'b00000000};
    rom_data[369]={8'b00010011,8'b00110000,8'b00000000};
    rom_data[373]={8'b00010011,8'b00101111,8'b00000000};
    rom_data[377]={8'b00010011,8'b00101110,8'b00000000};
    rom_data[381]={8'b00010011,8'b00101101,8'b00000000};
    rom_data[385]={8'b00010011,8'b00101100,8'b00000000};
    rom_data[389]={8'b00010011,8'b00101011,8'b00000000};
    rom_data[393]={8'b00010011,8'b00101010,8'b00000000};
    rom_data[397]={8'b00010011,8'b00101001,8'b00000000};
    rom_data[401]={8'b00010011,8'b00101000,8'b00000000};
    rom_data[405]={8'b00010011,8'b00100111,8'b00000000};
    rom_data[409]={8'b00010011,8'b00100110,8'b00000000};
    rom_data[413]={8'b00010011,8'b00100101,8'b00000000};
    rom_data[417]={8'b00010011,8'b00100100,8'b00000000};
    rom_data[421]={8'b00010011,8'b00100011,8'b00000000};
    rom_data[425]={8'b00010011,8'b00100010,8'b00000000};
    rom_data[429]={8'b00010011,8'b00100001,8'b00000000};
    rom_data[433]={8'b00010011,8'b00100000,8'b00000000};
    rom_data[437]={8'b00010011,8'b00011111,8'b00000000};
    rom_data[441]={8'b00010011,8'b00011110,8'b00000000};
    rom_data[445]={8'b00010011,8'b00011101,8'b00000000};
    rom_data[449]={8'b00010011,8'b00011100,8'b00000000};
    rom_data[453]={8'b00010011,8'b00011011,8'b00000000};
    rom_data[457]={8'b00010011,8'b00011010,8'b00000000};
    rom_data[461]={8'b00010011,8'b00011001,8'b00000000};
    rom_data[465]={8'b00010011,8'b00011000,8'b00000000};
    rom_data[469]={8'b00010011,8'b00010111,8'b00000000};
    rom_data[473]={8'b00010011,8'b00010110,8'b00000000};
    rom_data[477]={8'b00010011,8'b00010101,8'b00000000};
    rom_data[481]={8'b00010011,8'b00010100,8'b00000000};

    data_d = rom_data[addr];
  end
 

  always @(posedge clk) begin
    data_q <= data_d;
  end
 
endmodule