module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] addr,
    input go_home,
    // OUTPUT
    output [23:0] data,
    output rom_scan_is_done

  );
  
parameter rom_size = 641;

reg [15:0] rom_data [rom_size:0];
reg [23:0] data_d, data_q;
wire[14:0] addrs;
reg [15:0] antidata;
reg done;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;


reg [15:0] CH_A_d, CH_A_q;
reg [15:0] CH_B_d, CH_B_q;
reg [15:0] CH_C_d, CH_C_q;
reg [15:0] CH_D_d, CH_D_q;


assign data = data_q;
assign rom_scan_is_done = done;
assign addrs = addr[15:2];


always @(rst,addrs) begin
  if (rst) begin
      done = 1'b0;
  end else begin
      if (addrs == rom_size)
          done = 1'b1;
      else
          done = 1'b0;
  end     
end // always
 

always @(addrs) begin
    
    CH_A_d=CH_A_q;
    CH_B_d=CH_B_q;
    CH_C_d=CH_C_q;
    CH_D_d=CH_D_q;

    if (go_home==1'b1) begin
        case (addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (CH_A_q>home_bias) begin
                    CH_A_d=CH_A_q-home_step;
                end else if (CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_A_d=CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (CH_C_q>home_bias) begin
                    CH_C_d=CH_C_q-home_step;
                end else if (CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_C_d=CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (CH_B_q>home_bias) begin
                    CH_B_d=CH_B_q-home_step;
                end else if (CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_B_d=CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (CH_D_q>home_bias) begin
                    CH_D_d=CH_D_q-home_step;
                end else if (CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    CH_D_d=CH_D_q+home_step; 
                end 
            end

            default: begin
            end
        endcase

    end else begin // if go home==0
        case (addr[2:1])
            2'b00: begin
                CH_A_d= rom_data[addrs];
            end
            2'b01: begin
                CH_C_d= antidata;
            end
            2'b10: begin
                CH_B_d= rom_data[addrs];
            end
            2'b11: begin
                CH_D_d= antidata;
            end

        default: begin
            end
        endcase

    end // if go home 
end // always





always @(*) begin

  antidata = 16'hB900 - rom_data[addrs];


  rom_data[ 2]=16'b0010001010101010;
  rom_data[ 3]=16'b0101110110011100;
    rom_data[ 4]=16'b0010001010101010;
    rom_data[ 5]=16'b0110001110010101;
    rom_data[ 6]=16'b0010001100001010;
    rom_data[ 7]=16'b0110100101111100;
    rom_data[ 8]=16'b0010001110010000;
    rom_data[ 9]=16'b0110111101000100;
    rom_data[10]=16'b0010010000101001;
    rom_data[11]=16'b0111010011011101;
    rom_data[12]=16'b0010010011001110;
    rom_data[13]=16'b0111101000111010;
    rom_data[14]=16'b0010010101111001;
    rom_data[15]=16'b0111111101001110;
    rom_data[16]=16'b0010011000101001;
    rom_data[17]=16'b1000010000001100;
    rom_data[18]=16'b0010011011011011;
    rom_data[19]=16'b1000100001101001;
    rom_data[20]=16'b0010011110010001;
    rom_data[21]=16'b1000110001011001;
    rom_data[22]=16'b0010100001001000;
    rom_data[23]=16'b1000111111010100;
    rom_data[24]=16'b0010100100000000;
    rom_data[25]=16'b1001001011010000;
    rom_data[26]=16'b0010100110111001;
    rom_data[27]=16'b1001010101000110;
    rom_data[28]=16'b0010101001110100;
    rom_data[29]=16'b1001011100101111;
    rom_data[30]=16'b0010101100101111;
    rom_data[31]=16'b1001100010001001;
    rom_data[32]=16'b0010101111101010;
    rom_data[33]=16'b1001100101001110;
    rom_data[34]=16'b0010110010100110;
    rom_data[35]=16'b1001100101111101;
    rom_data[36]=16'b0010110101100010;
    rom_data[37]=16'b1001100100010110;
    rom_data[38]=16'b0010111000011111;
    rom_data[39]=16'b1001100000011010;
    rom_data[40]=16'b0010111011011100;
    rom_data[41]=16'b1001011010001011;
    rom_data[42]=16'b0010111110011001;
    rom_data[43]=16'b1001010001101100;
    rom_data[44]=16'b0011000001010110;
    rom_data[45]=16'b1001000111000100;
    rom_data[46]=16'b0011000100010100;
    rom_data[47]=16'b1000111010011000;
    rom_data[48]=16'b0011000111010010;
    rom_data[49]=16'b1000101011110001;
    rom_data[50]=16'b0011001010010000;
    rom_data[51]=16'b1000011011011000;
    rom_data[52]=16'b0011001101001110;
    rom_data[53]=16'b1000001001010110;
    rom_data[54]=16'b0011010000001100;
    rom_data[55]=16'b0111110101110110;
    rom_data[56]=16'b0011010011001010;
    rom_data[57]=16'b0111100001000110;
    rom_data[58]=16'b0011010110001000;
    rom_data[59]=16'b0111001011010001;
    rom_data[60]=16'b0011011001000111;
    rom_data[61]=16'b0110110100100101;
    rom_data[62]=16'b0011011100000101;
    rom_data[63]=16'b0110011101010000;
    rom_data[64]=16'b0011011111000100;
    rom_data[65]=16'b0110000101100000;
    rom_data[66]=16'b0011100010000010;
    rom_data[67]=16'b0101101101100100;
    rom_data[68]=16'b0011100101000001;
    rom_data[69]=16'b0101010101101011;
    rom_data[70]=16'b0011101000000000;
    rom_data[71]=16'b0100111110000100;
    rom_data[72]=16'b0011101010111110;
    rom_data[73]=16'b0100100110111100;
    rom_data[74]=16'b0011101101111101;
    rom_data[75]=16'b0100010000100011;
    rom_data[76]=16'b0011110000111100;
    rom_data[77]=16'b0011111011000110;
    rom_data[78]=16'b0011110011111011;
    rom_data[79]=16'b0011100110110010;
    rom_data[80]=16'b0011110110111001;
    rom_data[81]=16'b0011010011110100;
    rom_data[82]=16'b0011111001111000;
    rom_data[83]=16'b0011000010010111;
    rom_data[84]=16'b0011111100110111;
    rom_data[85]=16'b0010110010100111;
    rom_data[86]=16'b0011111111110110;
    rom_data[87]=16'b0010100100101100;
    rom_data[88]=16'b0100000010110101;
    rom_data[89]=16'b0010011000110000;
    rom_data[90]=16'b0100000101110100;
    rom_data[91]=16'b0010001110111010;
    rom_data[92]=16'b0100001000110011;
    rom_data[93]=16'b0010000111010001;
    rom_data[94]=16'b0100001011110010;
    rom_data[95]=16'b0010000001110111;
    rom_data[96]=16'b0100001110110001;
    rom_data[97]=16'b0001111110110010;
    rom_data[98]=16'b0100010001110000;
    rom_data[99]=16'b0001111110000011;
    rom_data[100]=16'b0100010100101111;
    rom_data[101]=16'b0001111111101010;
    rom_data[102]=16'b0100010111101110;
    rom_data[103]=16'b0010000011100110;
    rom_data[104]=16'b0100011010101101;
    rom_data[105]=16'b0010001001110101;
    rom_data[106]=16'b0100011101101100;
    rom_data[107]=16'b0010010010010100;
    rom_data[108]=16'b0100100000101011;
    rom_data[109]=16'b0010011100111100;
    rom_data[110]=16'b0100100011101010;
    rom_data[111]=16'b0010101001101000;
    rom_data[112]=16'b0100100110101001;
    rom_data[113]=16'b0010111000001111;
    rom_data[114]=16'b0100101001101000;
    rom_data[115]=16'b0011001000101000;
    rom_data[116]=16'b0100101100100111;
    rom_data[117]=16'b0011011010101010;
    rom_data[118]=16'b0100101111100110;
    rom_data[119]=16'b0011101110001010;
    rom_data[120]=16'b0100110010100101;
    rom_data[121]=16'b0100000010111010;
    rom_data[122]=16'b0100110101100100;
    rom_data[123]=16'b0100011000101111;
    rom_data[124]=16'b0100111000100011;
    rom_data[125]=16'b0100101111011011;
    rom_data[126]=16'b0100111011100001;
    rom_data[127]=16'b0101000110110000;
    rom_data[128]=16'b0100111110100000;
    rom_data[129]=16'b0101011110100000;
    rom_data[130]=16'b0101000001011111;
    rom_data[131]=16'b0101110110011100;
    rom_data[132]=16'b0101000100011110;
    rom_data[133]=16'b0110001110010101;
    rom_data[134]=16'b0101000111011101;
    rom_data[135]=16'b0110100101111100;
    rom_data[136]=16'b0101001010011100;
    rom_data[137]=16'b0110111101000100;
    rom_data[138]=16'b0101001101011011;
    rom_data[139]=16'b0111010011011101;
    rom_data[140]=16'b0101010000011010;
    rom_data[141]=16'b0111101000111010;
    rom_data[142]=16'b0101010011011001;
    rom_data[143]=16'b0111111101001110;
    rom_data[144]=16'b0101010110010111;
    rom_data[145]=16'b1000010000001100;
    rom_data[146]=16'b0101011001010110;
    rom_data[147]=16'b1000100001101001;
    rom_data[148]=16'b0101011100010101;
    rom_data[149]=16'b1000110001011001;
    rom_data[150]=16'b0101011111010100;
    rom_data[151]=16'b1000111111010100;
    rom_data[152]=16'b0101100010010011;
    rom_data[153]=16'b1001001011010000;
    rom_data[154]=16'b0101100101010001;
    rom_data[155]=16'b1001010101000110;
    rom_data[156]=16'b0101101000010000;
    rom_data[157]=16'b1001011100101111;
    rom_data[158]=16'b0101101011001111;
    rom_data[159]=16'b1001100010001001;
    rom_data[160]=16'b0101101110001101;
    rom_data[161]=16'b1001100101001110;
    rom_data[162]=16'b0101110001001100;
    rom_data[163]=16'b1001100101111101;
    rom_data[164]=16'b0101110100001011;
    rom_data[165]=16'b1001100100010110;
    rom_data[166]=16'b0101110111001001;
    rom_data[167]=16'b1001100000011010;
    rom_data[168]=16'b0101111010001000;
    rom_data[169]=16'b1001011010001011;
    rom_data[170]=16'b0101111101000110;
    rom_data[171]=16'b1001010001101100;
    rom_data[172]=16'b0110000000000101;
    rom_data[173]=16'b1001000111000100;
    rom_data[174]=16'b0110000011000011;
    rom_data[175]=16'b1000111010011000;
    rom_data[176]=16'b0110000110000001;
    rom_data[177]=16'b1000101011110001;
    rom_data[178]=16'b0110001001000000;
    rom_data[179]=16'b1000011011011000;
    rom_data[180]=16'b0110001011111110;
    rom_data[181]=16'b1000001001010110;
    rom_data[182]=16'b0110001110111100;
    rom_data[183]=16'b0111110101110110;
    rom_data[184]=16'b0110010001111010;
    rom_data[185]=16'b0111100001000110;
    rom_data[186]=16'b0110010100111001;
    rom_data[187]=16'b0111001011010001;
    rom_data[188]=16'b0110010111110111;
    rom_data[189]=16'b0110110100100101;
    rom_data[190]=16'b0110011010110101;
    rom_data[191]=16'b0110011101010000;
    rom_data[192]=16'b0110011101110011;
    rom_data[193]=16'b0110000101100000;
    rom_data[194]=16'b0110100000110001;
    rom_data[195]=16'b0101101101100100;
    rom_data[196]=16'b0110100011101110;
    rom_data[197]=16'b0101010101101011;
    rom_data[198]=16'b0110100110101100;
    rom_data[199]=16'b0100111110000100;
    rom_data[200]=16'b0110101001101010;
    rom_data[201]=16'b0100100110111100;
    rom_data[202]=16'b0110101100101000;
    rom_data[203]=16'b0100010000100011;
    rom_data[204]=16'b0110101111100101;
    rom_data[205]=16'b0011111011000110;
    rom_data[206]=16'b0110110010100011;
    rom_data[207]=16'b0011100110110010;
    rom_data[208]=16'b0110110101100000;
    rom_data[209]=16'b0011010011110100;
    rom_data[210]=16'b0110111000011110;
    rom_data[211]=16'b0011000010010111;
    rom_data[212]=16'b0110111011011011;
    rom_data[213]=16'b0010110010100111;
    rom_data[214]=16'b0110111110011000;
    rom_data[215]=16'b0010100100101100;
    rom_data[216]=16'b0111000001010101;
    rom_data[217]=16'b0010011000110000;
    rom_data[218]=16'b0111000100010010;
    rom_data[219]=16'b0010001110111010;
    rom_data[220]=16'b0111000111001111;
    rom_data[221]=16'b0010000111010001;
    rom_data[222]=16'b0111001010001011;
    rom_data[223]=16'b0010000001110111;
    rom_data[224]=16'b0111001101001000;
    rom_data[225]=16'b0001111110110010;
    rom_data[226]=16'b0111010000000100;
    rom_data[227]=16'b0001111110000011;
    rom_data[228]=16'b0111010011000001;
    rom_data[229]=16'b0001111111101010;
    rom_data[230]=16'b0111010101111101;
    rom_data[231]=16'b0010000011100110;
    rom_data[232]=16'b0111011000111001;
    rom_data[233]=16'b0010001001110101;
    rom_data[234]=16'b0111011011110101;
    rom_data[235]=16'b0010010010010100;
    rom_data[236]=16'b0111011110110000;
    rom_data[237]=16'b0010011100111100;
    rom_data[238]=16'b0111100001101100;
    rom_data[239]=16'b0010101001101000;
    rom_data[240]=16'b0111100100100111;
    rom_data[241]=16'b0010111000001111;
    rom_data[242]=16'b0111100111100010;
    rom_data[243]=16'b0011001000101000;
    rom_data[244]=16'b0111101010011101;
    rom_data[245]=16'b0011011010101010;
    rom_data[246]=16'b0111101101011000;
    rom_data[247]=16'b0011101110001010;
    rom_data[248]=16'b0111110000010010;
    rom_data[249]=16'b0100000010111010;
    rom_data[250]=16'b0111110011001100;
    rom_data[251]=16'b0100011000101111;
    rom_data[252]=16'b0111110110000110;
    rom_data[253]=16'b0100101111011011;
    rom_data[254]=16'b0111111001000000;
    rom_data[255]=16'b0101000110110000;
    rom_data[256]=16'b0111111011111001;
    rom_data[257]=16'b0101011110100000;
    rom_data[258]=16'b0111111110110010;
    rom_data[259]=16'b0101110110011100;
    rom_data[260]=16'b1000000001101011;
    rom_data[261]=16'b0110001110010101;
    rom_data[262]=16'b1000000100100011;
    rom_data[263]=16'b0110100101111100;
    rom_data[264]=16'b1000000111011011;
    rom_data[265]=16'b0110111101000100;
    rom_data[266]=16'b1000001010010010;
    rom_data[267]=16'b0111010011011101;
    rom_data[268]=16'b1000001101001001;
    rom_data[269]=16'b0111101000111010;
    rom_data[270]=16'b1000001111111111;
    rom_data[271]=16'b0111111101001110;
    rom_data[272]=16'b1000010010110101;
    rom_data[273]=16'b1000010000001100;
    rom_data[274]=16'b1000010101101010;
    rom_data[275]=16'b1000100001101001;
    rom_data[276]=16'b1000011000011111;
    rom_data[277]=16'b1000110001011001;
    rom_data[278]=16'b1000011011010011;
    rom_data[279]=16'b1000111111010100;
    rom_data[280]=16'b1000011110000110;
    rom_data[281]=16'b1001001011010000;
    rom_data[282]=16'b1000100000111000;
    rom_data[283]=16'b1001010101000110;
    rom_data[284]=16'b1000100011101001;
    rom_data[285]=16'b1001011100101111;
    rom_data[286]=16'b1000100110011010;
    rom_data[287]=16'b1001100010001001;
    rom_data[288]=16'b1000101001001001;
    rom_data[289]=16'b1001100101001110;
    rom_data[290]=16'b1000101011111000;
    rom_data[291]=16'b1001100101111101;
    rom_data[292]=16'b1000101110100101;
    rom_data[293]=16'b1001100100010110;
    rom_data[294]=16'b1000110001010000;
    rom_data[295]=16'b1001100000011010;
    rom_data[296]=16'b1000110011111010;
    rom_data[297]=16'b1001011010001011;
    rom_data[298]=16'b1000110110100011;
    rom_data[299]=16'b1001010001101100;
    rom_data[300]=16'b1000111001001001;
    rom_data[301]=16'b1001000111000100;
    rom_data[302]=16'b1000111011101110;
    rom_data[303]=16'b1000111010011000;
    rom_data[304]=16'b1000111110010000;
    rom_data[305]=16'b1000101011110001;
    rom_data[306]=16'b1001000000110000;
    rom_data[307]=16'b1000011011011000;
    rom_data[308]=16'b1001000011001101;
    rom_data[309]=16'b1000001001010110;
    rom_data[310]=16'b1001000101100111;
    rom_data[311]=16'b0111110101110110;
    rom_data[312]=16'b1001000111111101;
    rom_data[313]=16'b0111100001000110;
    rom_data[314]=16'b1001001010010000;
    rom_data[315]=16'b0111001011010001;
    rom_data[316]=16'b1001001100011110;
    rom_data[317]=16'b0110110100100101;
    rom_data[318]=16'b1001001110100110;
    rom_data[319]=16'b0110011101010000;
    rom_data[320]=16'b1001010000101001;
    rom_data[321]=16'b0110000101100000;
    rom_data[322]=16'b1001010000101001;
    rom_data[323]=16'b0101101101100100;
    rom_data[324]=16'b1001001110100110;
    rom_data[325]=16'b0101010101101011;
    rom_data[326]=16'b1001001100011110;
    rom_data[327]=16'b0100111110000100;
    rom_data[328]=16'b1001001010010000;
    rom_data[329]=16'b0100100110111100;
    rom_data[330]=16'b1001000111111101;
    rom_data[331]=16'b0100010000100011;
    rom_data[332]=16'b1001000101100111;
    rom_data[333]=16'b0011111011000110;
    rom_data[334]=16'b1001000011001101;
    rom_data[335]=16'b0011100110110010;
    rom_data[336]=16'b1001000000110000;
    rom_data[337]=16'b0011010011110100;
    rom_data[338]=16'b1000111110010000;
    rom_data[339]=16'b0011000010010111;
    rom_data[340]=16'b1000111011101110;
    rom_data[341]=16'b0010110010100111;
    rom_data[342]=16'b1000111001001001;
    rom_data[343]=16'b0010100100101100;
    rom_data[344]=16'b1000110110100011;
    rom_data[345]=16'b0010011000110000;
    rom_data[346]=16'b1000110011111010;
    rom_data[347]=16'b0010001110111010;
    rom_data[348]=16'b1000110001010000;
    rom_data[349]=16'b0010000111010001;
    rom_data[350]=16'b1000101110100101;
    rom_data[351]=16'b0010000001110111;
    rom_data[352]=16'b1000101011111000;
    rom_data[353]=16'b0001111110110010;
    rom_data[354]=16'b1000101001001001;
    rom_data[355]=16'b0001111110000011;
    rom_data[356]=16'b1000100110011010;
    rom_data[357]=16'b0001111111101010;
    rom_data[358]=16'b1000100011101001;
    rom_data[359]=16'b0010000011100110;
    rom_data[360]=16'b1000100000111000;
    rom_data[361]=16'b0010001001110101;
    rom_data[362]=16'b1000011110000110;
    rom_data[363]=16'b0010010010010100;
    rom_data[364]=16'b1000011011010011;
    rom_data[365]=16'b0010011100111100;
    rom_data[366]=16'b1000011000011111;
    rom_data[367]=16'b0010101001101000;
    rom_data[368]=16'b1000010101101010;
    rom_data[369]=16'b0010111000001111;
    rom_data[370]=16'b1000010010110101;
    rom_data[371]=16'b0011001000101000;
    rom_data[372]=16'b1000001111111111;
    rom_data[373]=16'b0011011010101010;
    rom_data[374]=16'b1000001101001001;
    rom_data[375]=16'b0011101110001010;
    rom_data[376]=16'b1000001010010010;
    rom_data[377]=16'b0100000010111010;
    rom_data[378]=16'b1000000111011011;
    rom_data[379]=16'b0100011000101111;
    rom_data[380]=16'b1000000100100011;
    rom_data[381]=16'b0100101111011011;
    rom_data[382]=16'b1000000001101011;
    rom_data[383]=16'b0101000110110000;
    rom_data[384]=16'b0111111110110010;
    rom_data[385]=16'b0101011110100000;
    rom_data[386]=16'b0111111011111001;
    rom_data[387]=16'b0101110110011100;
    rom_data[388]=16'b0111111001000000;
    rom_data[389]=16'b0110001110010101;
    rom_data[390]=16'b0111110110000110;
    rom_data[391]=16'b0110100101111100;
    rom_data[392]=16'b0111110011001100;
    rom_data[393]=16'b0110111101000100;
    rom_data[394]=16'b0111110000010010;
    rom_data[395]=16'b0111010011011101;
    rom_data[396]=16'b0111101101011000;
    rom_data[397]=16'b0111101000111010;
    rom_data[398]=16'b0111101010011101;
    rom_data[399]=16'b0111111101001110;
    rom_data[400]=16'b0111100111100010;
    rom_data[401]=16'b1000010000001100;
    rom_data[402]=16'b0111100100100111;
    rom_data[403]=16'b1000100001101001;
    rom_data[404]=16'b0111100001101100;
    rom_data[405]=16'b1000110001011001;
    rom_data[406]=16'b0111011110110000;
    rom_data[407]=16'b1000111111010100;
    rom_data[408]=16'b0111011011110101;
    rom_data[409]=16'b1001001011010000;
    rom_data[410]=16'b0111011000111001;
    rom_data[411]=16'b1001010101000110;
    rom_data[412]=16'b0111010101111101;
    rom_data[413]=16'b1001011100101111;
    rom_data[414]=16'b0111010011000001;
    rom_data[415]=16'b1001100010001001;
    rom_data[416]=16'b0111010000000100;
    rom_data[417]=16'b1001100101001110;
    rom_data[418]=16'b0111001101001000;
    rom_data[419]=16'b1001100101111101;
    rom_data[420]=16'b0111001010001011;
    rom_data[421]=16'b1001100100010110;
    rom_data[422]=16'b0111000111001111;
    rom_data[423]=16'b1001100000011010;
    rom_data[424]=16'b0111000100010010;
    rom_data[425]=16'b1001011010001011;
    rom_data[426]=16'b0111000001010101;
    rom_data[427]=16'b1001010001101100;
    rom_data[428]=16'b0110111110011000;
    rom_data[429]=16'b1001000111000100;
    rom_data[430]=16'b0110111011011011;
    rom_data[431]=16'b1000111010011000;
    rom_data[432]=16'b0110111000011110;
    rom_data[433]=16'b1000101011110001;
    rom_data[434]=16'b0110110101100000;
    rom_data[435]=16'b1000011011011000;
    rom_data[436]=16'b0110110010100011;
    rom_data[437]=16'b1000001001010110;
    rom_data[438]=16'b0110101111100101;
    rom_data[439]=16'b0111110101110110;
    rom_data[440]=16'b0110101100101000;
    rom_data[441]=16'b0111100001000110;
    rom_data[442]=16'b0110101001101010;
    rom_data[443]=16'b0111001011010001;
    rom_data[444]=16'b0110100110101100;
    rom_data[445]=16'b0110110100100101;
    rom_data[446]=16'b0110100011101110;
    rom_data[447]=16'b0110011101010000;
    rom_data[448]=16'b0110100000110001;
    rom_data[449]=16'b0110000101100000;
    rom_data[450]=16'b0110011101110011;
    rom_data[451]=16'b0101101101100100;
    rom_data[452]=16'b0110011010110101;
    rom_data[453]=16'b0101010101101011;
    rom_data[454]=16'b0110010111110111;
    rom_data[455]=16'b0100111110000100;
    rom_data[456]=16'b0110010100111001;
    rom_data[457]=16'b0100100110111100;
    rom_data[458]=16'b0110010001111010;
    rom_data[459]=16'b0100010000100011;
    rom_data[460]=16'b0110001110111100;
    rom_data[461]=16'b0011111011000110;
    rom_data[462]=16'b0110001011111110;
    rom_data[463]=16'b0011100110110010;
    rom_data[464]=16'b0110001001000000;
    rom_data[465]=16'b0011010011110100;
    rom_data[466]=16'b0110000110000001;
    rom_data[467]=16'b0011000010010111;
    rom_data[468]=16'b0110000011000011;
    rom_data[469]=16'b0010110010100111;
    rom_data[470]=16'b0110000000000101;
    rom_data[471]=16'b0010100100101100;
    rom_data[472]=16'b0101111101000110;
    rom_data[473]=16'b0010011000110000;
    rom_data[474]=16'b0101111010001000;
    rom_data[475]=16'b0010001110111010;
    rom_data[476]=16'b0101110111001001;
    rom_data[477]=16'b0010000111010001;
    rom_data[478]=16'b0101110100001011;
    rom_data[479]=16'b0010000001110111;
    rom_data[480]=16'b0101110001001100;
    rom_data[481]=16'b0001111110110010;
    rom_data[482]=16'b0101101110001101;
    rom_data[483]=16'b0001111110000011;
    rom_data[484]=16'b0101101011001111;
    rom_data[485]=16'b0001111111101010;
    rom_data[486]=16'b0101101000010000;
    rom_data[487]=16'b0010000011100110;
    rom_data[488]=16'b0101100101010001;
    rom_data[489]=16'b0010001001110101;
    rom_data[490]=16'b0101100010010011;
    rom_data[491]=16'b0010010010010100;
    rom_data[492]=16'b0101011111010100;
    rom_data[493]=16'b0010011100111100;
    rom_data[494]=16'b0101011100010101;
    rom_data[495]=16'b0010101001101000;
    rom_data[496]=16'b0101011001010110;
    rom_data[497]=16'b0010111000001111;
    rom_data[498]=16'b0101010110010111;
    rom_data[499]=16'b0011001000101000;
    rom_data[500]=16'b0101010011011001;
    rom_data[501]=16'b0011011010101010;
    rom_data[502]=16'b0101010000011010;
    rom_data[503]=16'b0011101110001010;
    rom_data[504]=16'b0101001101011011;
    rom_data[505]=16'b0100000010111010;
    rom_data[506]=16'b0101001010011100;
    rom_data[507]=16'b0100011000101111;
    rom_data[508]=16'b0101000111011101;
    rom_data[509]=16'b0100101111011011;
    rom_data[510]=16'b0101000100011110;
    rom_data[511]=16'b0101000110110000;
    rom_data[512]=16'b0101000001011111;
    rom_data[513]=16'b0101011110100000;
    rom_data[514]=16'b0100111110100000;
    rom_data[515]=16'b0101110110011100;
    rom_data[516]=16'b0100111011100001;
    rom_data[517]=16'b0110001110010101;
    rom_data[518]=16'b0100111000100011;
    rom_data[519]=16'b0110100101111100;
    rom_data[520]=16'b0100110101100100;
    rom_data[521]=16'b0110111101000100;
    rom_data[522]=16'b0100110010100101;
    rom_data[523]=16'b0111010011011101;
    rom_data[524]=16'b0100101111100110;
    rom_data[525]=16'b0111101000111010;
    rom_data[526]=16'b0100101100100111;
    rom_data[527]=16'b0111111101001110;
    rom_data[528]=16'b0100101001101000;
    rom_data[529]=16'b1000010000001100;
    rom_data[530]=16'b0100100110101001;
    rom_data[531]=16'b1000100001101001;
    rom_data[532]=16'b0100100011101010;
    rom_data[533]=16'b1000110001011001;
    rom_data[534]=16'b0100100000101011;
    rom_data[535]=16'b1000111111010100;
    rom_data[536]=16'b0100011101101100;
    rom_data[537]=16'b1001001011010000;
    rom_data[538]=16'b0100011010101101;
    rom_data[539]=16'b1001010101000110;
    rom_data[540]=16'b0100010111101110;
    rom_data[541]=16'b1001011100101111;
    rom_data[542]=16'b0100010100101111;
    rom_data[543]=16'b1001100010001001;
    rom_data[544]=16'b0100010001110000;
    rom_data[545]=16'b1001100101001110;
    rom_data[546]=16'b0100001110110001;
    rom_data[547]=16'b1001100101111101;
    rom_data[548]=16'b0100001011110010;
    rom_data[549]=16'b1001100100010110;
    rom_data[550]=16'b0100001000110011;
    rom_data[551]=16'b1001100000011010;
    rom_data[552]=16'b0100000101110100;
    rom_data[553]=16'b1001011010001011;
    rom_data[554]=16'b0100000010110101;
    rom_data[555]=16'b1001010001101100;
    rom_data[556]=16'b0011111111110110;
    rom_data[557]=16'b1001000111000100;
    rom_data[558]=16'b0011111100110111;
    rom_data[559]=16'b1000111010011000;
    rom_data[560]=16'b0011111001111000;
    rom_data[561]=16'b1000101011110001;
    rom_data[562]=16'b0011110110111001;
    rom_data[563]=16'b1000011011011000;
    rom_data[564]=16'b0011110011111011;
    rom_data[565]=16'b1000001001010110;
    rom_data[566]=16'b0011110000111100;
    rom_data[567]=16'b0111110101110110;
    rom_data[568]=16'b0011101101111101;
    rom_data[569]=16'b0111100001000110;
    rom_data[570]=16'b0011101010111110;
    rom_data[571]=16'b0111001011010001;
    rom_data[572]=16'b0011101000000000;
    rom_data[573]=16'b0110110100100101;
    rom_data[574]=16'b0011100101000001;
    rom_data[575]=16'b0110011101010000;
    rom_data[576]=16'b0011100010000010;
    rom_data[577]=16'b0110000101100000;
    rom_data[578]=16'b0011011111000100;
    rom_data[579]=16'b0101101101100100;
    rom_data[580]=16'b0011011100000101;
    rom_data[581]=16'b0101010101101011;
    rom_data[582]=16'b0011011001000111;
    rom_data[583]=16'b0100111110000100;
    rom_data[584]=16'b0011010110001000;
    rom_data[585]=16'b0100100110111100;
    rom_data[586]=16'b0011010011001010;
    rom_data[587]=16'b0100010000100011;
    rom_data[588]=16'b0011010000001100;
    rom_data[589]=16'b0011111011000110;
    rom_data[590]=16'b0011001101001110;
    rom_data[591]=16'b0011100110110010;
    rom_data[592]=16'b0011001010010000;
    rom_data[593]=16'b0011010011110100;
    rom_data[594]=16'b0011000111010010;
    rom_data[595]=16'b0011000010010111;
    rom_data[596]=16'b0011000100010100;
    rom_data[597]=16'b0010110010100111;
    rom_data[598]=16'b0011000001010110;
    rom_data[599]=16'b0010100100101100;
    rom_data[600]=16'b0010111110011001;
    rom_data[601]=16'b0010011000110000;
    rom_data[602]=16'b0010111011011100;
    rom_data[603]=16'b0010001110111010;
    rom_data[604]=16'b0010111000011111;
    rom_data[605]=16'b0010000111010001;
    rom_data[606]=16'b0010110101100010;
    rom_data[607]=16'b0010000001110111;
    rom_data[608]=16'b0010110010100110;
    rom_data[609]=16'b0001111110110010;
    rom_data[610]=16'b0010101111101010;
    rom_data[611]=16'b0001111110000011;
    rom_data[612]=16'b0010101100101111;
    rom_data[613]=16'b0001111111101010;
    rom_data[614]=16'b0010101001110100;
    rom_data[615]=16'b0010000011100110;
    rom_data[616]=16'b0010100110111001;
    rom_data[617]=16'b0010001001110101;
    rom_data[618]=16'b0010100100000000;
    rom_data[619]=16'b0010010010010100;
    rom_data[620]=16'b0010100001001000;
    rom_data[621]=16'b0010011100111100;
    rom_data[622]=16'b0010011110010001;
    rom_data[623]=16'b0010101001101000;
    rom_data[624]=16'b0010011011011011;
    rom_data[625]=16'b0010111000001111;
    rom_data[626]=16'b0010011000101001;
    rom_data[627]=16'b0011001000101000;
    rom_data[628]=16'b0010010101111001;
    rom_data[629]=16'b0011011010101010;
    rom_data[630]=16'b0010010011001110;
    rom_data[631]=16'b0011101110001010;
    rom_data[632]=16'b0010010000101001;
    rom_data[633]=16'b0100000010111010;
    rom_data[634]=16'b0010001110010000;
    rom_data[635]=16'b0100011000101111;
    rom_data[636]=16'b0010001100001010;
    rom_data[637]=16'b0100101111011011;
    rom_data[638]=16'b0010001010101010;
    rom_data[639]=16'b0101000110110000;
    rom_data[640]=16'b0010001010101010;
    rom_data[641]=16'b0101011110100000;





    if (addr[0]==1'b0) begin
        data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
    end else begin //data in 50%
        
        case (addr[2:1])
            2'b00: begin // this is a CHANNEL A
                data_d = {6'b000110, addr[2:1], CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                data_d = {6'b000110, addr[2:1], CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                data_d = {6'b000110, addr[2:1], CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                data_d = {6'b000110, addr[2:1], CH_D_q};
            end

            default: begin
            end
        endcase

    end // if VREF
end // always


always @(posedge addr[0]) begin
    CH_A_q<=CH_A_d;
    CH_B_q<=CH_B_d;
    CH_C_q<=CH_C_d;
    CH_D_q<=CH_D_d;
end


always @(posedge clk) begin
  if (addr==0) begin
    data_q <= 24'b001010000000000000000001; // SOFT_RESET;//
  end else if (addr==1) begin
    data_q <= 24'b00111000_0000000000000000;    //Vref 
  end else begin
    data_q <= data_d;
  end
end // always
 
endmodule