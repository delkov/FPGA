 39 lines, assign
 
module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] f1_addr,
    input [15:0] f2_addr,
    input [15:0] f3_addr,
    input [15:0] f4_addr,
    input [15:0] f5_addr,
    input [15:0] f6_addr,

    input go_home,
    // OUTPUT
    output [23:0] f1_data,
    output [23:0] f2_data,
    output [23:0] f3_data,
    output [23:0] f4_data,
    output [23:0] f5_data,
    output [23:0] f6_data
  );
  
parameter rom_size = 14041;

wire [7:0] rom_data [rom_size:0];

   assign rom_data[ 2]=8'b00101100;
   assign rom_data[ 3]=8'b01011011;
   assign rom_data[ 4]=8'b00101100;
   assign rom_data[ 5]=8'b01011100;
   assign rom_data[ 6]=8'b00101100;
   assign rom_data[ 7]=8'b01011110;
   assign rom_data[ 8]=8'b00101100;
   assign rom_data[ 9]=8'b01011111;
   assign rom_data[10]=8'b00101100;
   assign rom_data[11]=8'b01100001;
   assign rom_data[12]=8'b00101100;
   assign rom_data[13]=8'b01100010;
   assign rom_data[14]=8'b00101100;
   assign rom_data[15]=8'b01100011;
   assign rom_data[16]=8'b00101100;
   assign rom_data[17]=8'b01100101;
   assign rom_data[18]=8'b00101100;
   assign rom_data[19]=8'b01100110;
   assign rom_data[20]=8'b00101100;
   assign rom_data[21]=8'b01100111;
   assign rom_data[22]=8'b00101100;
   assign rom_data[23]=8'b01101001;
   assign rom_data[24]=8'b00101100;
   assign rom_data[25]=8'b01101010;
   assign rom_data[26]=8'b00101100;
   assign rom_data[27]=8'b01101100;
   assign rom_data[28]=8'b00101100;
   assign rom_data[29]=8'b01101101;
   assign rom_data[30]=8'b00101100;
   assign rom_data[31]=8'b01101110;
   assign rom_data[32]=8'b00101100;
   assign rom_data[33]=8'b01110000;
   assign rom_data[34]=8'b00101101;
   assign rom_data[35]=8'b01110001;
   assign rom_data[36]=8'b00101101;
   assign rom_data[37]=8'b01110010;
   assign rom_data[38]=8'b00101101;
   assign rom_data[39]=8'b01110100;
   assign rom_data[40]=8'b00101101;
   assign rom_data[41]=8'b01110101;
   assign rom_data[42]=8'b00101101;
   assign rom_data[43]=8'b01110110;
   assign rom_data[44]=8'b00101101;
   assign rom_data[45]=8'b01110111;
   assign rom_data[46]=8'b00101101;
   assign rom_data[47]=8'b01111001;
   assign rom_data[48]=8'b00101101;
   assign rom_data[49]=8'b01111010;
   assign rom_data[50]=8'b00101101;
   assign rom_data[51]=8'b01111011;
   assign rom_data[52]=8'b00101101;
   assign rom_data[53]=8'b01111100;
   assign rom_data[54]=8'b00101101;
   assign rom_data[55]=8'b01111101;
   assign rom_data[56]=8'b00101101;
   assign rom_data[57]=8'b01111110;
   assign rom_data[58]=8'b00101101;
   assign rom_data[59]=8'b01111111;
   assign rom_data[60]=8'b00101101;
   assign rom_data[61]=8'b10000000;
   assign rom_data[62]=8'b00101101;
   assign rom_data[63]=8'b10000001;
   assign rom_data[64]=8'b00101101;
   assign rom_data[65]=8'b10000010;
   assign rom_data[66]=8'b00101101;
   assign rom_data[67]=8'b10000011;
   assign rom_data[68]=8'b00101101;
   assign rom_data[69]=8'b10000100;
   assign rom_data[70]=8'b00101101;
   assign rom_data[71]=8'b10000101;
   assign rom_data[72]=8'b00101101;
   assign rom_data[73]=8'b10000110;
   assign rom_data[74]=8'b00101101;
   assign rom_data[75]=8'b10000110;
   assign rom_data[76]=8'b00101101;
   assign rom_data[77]=8'b10000111;
   assign rom_data[78]=8'b00101101;
   assign rom_data[79]=8'b10001000;
   assign rom_data[80]=8'b00101101;
   assign rom_data[81]=8'b10001000;
   assign rom_data[82]=8'b00101101;
   assign rom_data[83]=8'b10001001;
   assign rom_data[84]=8'b00101101;
   assign rom_data[85]=8'b10001001;
   assign rom_data[86]=8'b00101101;
   assign rom_data[87]=8'b10001001;
   assign rom_data[88]=8'b00101101;
   assign rom_data[89]=8'b10001010;
   assign rom_data[90]=8'b00101101;
   assign rom_data[91]=8'b10001010;
   assign rom_data[92]=8'b00101101;
   assign rom_data[93]=8'b10001010;
   assign rom_data[94]=8'b00101101;
   assign rom_data[95]=8'b10001010;
   assign rom_data[96]=8'b00101101;
   assign rom_data[97]=8'b10001010;
   assign rom_data[98]=8'b00101101;
   assign rom_data[99]=8'b10001001;
   assign rom_data[100]=8'b00101101;
   assign rom_data[101]=8'b10001001;
   assign rom_data[102]=8'b00101101;
   assign rom_data[103]=8'b10001001;
   assign rom_data[104]=8'b00101101;
   assign rom_data[105]=8'b10001000;
   assign rom_data[106]=8'b00101101;
   assign rom_data[107]=8'b10001000;
   assign rom_data[108]=8'b00101101;
   assign rom_data[109]=8'b10000111;
   assign rom_data[110]=8'b00101110;
   assign rom_data[111]=8'b10000111;
   assign rom_data[112]=8'b00101110;
   assign rom_data[113]=8'b10000110;
   assign rom_data[114]=8'b00101110;
   assign rom_data[115]=8'b10000101;
   assign rom_data[116]=8'b00101110;
   assign rom_data[117]=8'b10000100;
   assign rom_data[118]=8'b00101110;
   assign rom_data[119]=8'b10000011;
   assign rom_data[120]=8'b00101110;
   assign rom_data[121]=8'b10000011;
   assign rom_data[122]=8'b00101110;
   assign rom_data[123]=8'b10000010;
   assign rom_data[124]=8'b00101110;
   assign rom_data[125]=8'b10000001;
   assign rom_data[126]=8'b00101110;
   assign rom_data[127]=8'b10000000;
   assign rom_data[128]=8'b00101110;
   assign rom_data[129]=8'b01111110;
   assign rom_data[130]=8'b00101110;
   assign rom_data[131]=8'b01111101;
   assign rom_data[132]=8'b00101110;
   assign rom_data[133]=8'b01111100;
   assign rom_data[134]=8'b00101110;
   assign rom_data[135]=8'b01111011;
   assign rom_data[136]=8'b00101110;
   assign rom_data[137]=8'b01111010;
   assign rom_data[138]=8'b00101110;
   assign rom_data[139]=8'b01111001;
   assign rom_data[140]=8'b00101110;
   assign rom_data[141]=8'b01110111;
   assign rom_data[142]=8'b00101110;
   assign rom_data[143]=8'b01110110;
   assign rom_data[144]=8'b00101110;
   assign rom_data[145]=8'b01110101;
   assign rom_data[146]=8'b00101110;
   assign rom_data[147]=8'b01110100;
   assign rom_data[148]=8'b00101110;
   assign rom_data[149]=8'b01110010;
   assign rom_data[150]=8'b00101110;
   assign rom_data[151]=8'b01110001;
   assign rom_data[152]=8'b00101110;
   assign rom_data[153]=8'b01110000;
   assign rom_data[154]=8'b00101110;
   assign rom_data[155]=8'b01101110;
   assign rom_data[156]=8'b00101110;
   assign rom_data[157]=8'b01101101;
   assign rom_data[158]=8'b00101110;
   assign rom_data[159]=8'b01101100;
   assign rom_data[160]=8'b00101110;
   assign rom_data[161]=8'b01101010;
   assign rom_data[162]=8'b00101110;
   assign rom_data[163]=8'b01101001;
   assign rom_data[164]=8'b00101110;
   assign rom_data[165]=8'b01101000;
   assign rom_data[166]=8'b00101110;
   assign rom_data[167]=8'b01100110;
   assign rom_data[168]=8'b00101110;
   assign rom_data[169]=8'b01100101;
   assign rom_data[170]=8'b00101110;
   assign rom_data[171]=8'b01100011;
   assign rom_data[172]=8'b00101110;
   assign rom_data[173]=8'b01100010;
   assign rom_data[174]=8'b00101110;
   assign rom_data[175]=8'b01100001;
   assign rom_data[176]=8'b00101110;
   assign rom_data[177]=8'b01011111;
   assign rom_data[178]=8'b00101110;
   assign rom_data[179]=8'b01011110;
   assign rom_data[180]=8'b00101110;
   assign rom_data[181]=8'b01011100;
   assign rom_data[182]=8'b00101110;
   assign rom_data[183]=8'b01011011;
   assign rom_data[184]=8'b00101110;
   assign rom_data[185]=8'b01011010;
   assign rom_data[186]=8'b00101110;
   assign rom_data[187]=8'b01011000;
   assign rom_data[188]=8'b00101111;
   assign rom_data[189]=8'b01010111;
   assign rom_data[190]=8'b00101111;
   assign rom_data[191]=8'b01010101;
   assign rom_data[192]=8'b00101111;
   assign rom_data[193]=8'b01010100;
   assign rom_data[194]=8'b00101111;
   assign rom_data[195]=8'b01010010;
   assign rom_data[196]=8'b00101111;
   assign rom_data[197]=8'b01010001;
   assign rom_data[198]=8'b00101111;
   assign rom_data[199]=8'b01010000;
   assign rom_data[200]=8'b00101111;
   assign rom_data[201]=8'b01001110;
   assign rom_data[202]=8'b00101111;
   assign rom_data[203]=8'b01001101;
   assign rom_data[204]=8'b00101111;
   assign rom_data[205]=8'b01001100;
   assign rom_data[206]=8'b00101111;
   assign rom_data[207]=8'b01001010;
   assign rom_data[208]=8'b00101111;
   assign rom_data[209]=8'b01001001;
   assign rom_data[210]=8'b00101111;
   assign rom_data[211]=8'b01001000;
   assign rom_data[212]=8'b00101111;
   assign rom_data[213]=8'b01000110;
   assign rom_data[214]=8'b00101111;
   assign rom_data[215]=8'b01000101;
   assign rom_data[216]=8'b00101111;
   assign rom_data[217]=8'b01000100;
   assign rom_data[218]=8'b00101111;
   assign rom_data[219]=8'b01000010;
   assign rom_data[220]=8'b00101111;
   assign rom_data[221]=8'b01000001;
   assign rom_data[222]=8'b00101111;
   assign rom_data[223]=8'b01000000;
   assign rom_data[224]=8'b00101111;
   assign rom_data[225]=8'b00111111;
   assign rom_data[226]=8'b00101111;
   assign rom_data[227]=8'b00111101;
   assign rom_data[228]=8'b00101111;
   assign rom_data[229]=8'b00111100;
   assign rom_data[230]=8'b00101111;
   assign rom_data[231]=8'b00111011;
   assign rom_data[232]=8'b00101111;
   assign rom_data[233]=8'b00111010;
   assign rom_data[234]=8'b00101111;
   assign rom_data[235]=8'b00111001;
   assign rom_data[236]=8'b00101111;
   assign rom_data[237]=8'b00111000;
   assign rom_data[238]=8'b00101111;
   assign rom_data[239]=8'b00110110;
   assign rom_data[240]=8'b00101111;
   assign rom_data[241]=8'b00110101;
   assign rom_data[242]=8'b00101111;
   assign rom_data[243]=8'b00110100;
   assign rom_data[244]=8'b00101111;
   assign rom_data[245]=8'b00110011;
   assign rom_data[246]=8'b00101111;
   assign rom_data[247]=8'b00110011;
   assign rom_data[248]=8'b00101111;
   assign rom_data[249]=8'b00110010;
   assign rom_data[250]=8'b00101111;
   assign rom_data[251]=8'b00110001;
   assign rom_data[252]=8'b00101111;
   assign rom_data[253]=8'b00110000;
   assign rom_data[254]=8'b00101111;
   assign rom_data[255]=8'b00101111;
   assign rom_data[256]=8'b00101111;
   assign rom_data[257]=8'b00101111;
   assign rom_data[258]=8'b00101111;
   assign rom_data[259]=8'b00101110;
   assign rom_data[260]=8'b00101111;
   assign rom_data[261]=8'b00101110;
   assign rom_data[262]=8'b00101111;
   assign rom_data[263]=8'b00101101;
   assign rom_data[264]=8'b00110000;
   assign rom_data[265]=8'b00101101;
   assign rom_data[266]=8'b00110000;
   assign rom_data[267]=8'b00101100;
   assign rom_data[268]=8'b00110000;
   assign rom_data[269]=8'b00101100;
   assign rom_data[270]=8'b00110000;
   assign rom_data[271]=8'b00101100;
   assign rom_data[272]=8'b00110000;
   assign rom_data[273]=8'b00101100;
   assign rom_data[274]=8'b00110000;
   assign rom_data[275]=8'b00101100;
   assign rom_data[276]=8'b00110000;
   assign rom_data[277]=8'b00101100;
   assign rom_data[278]=8'b00110000;
   assign rom_data[279]=8'b00101100;
   assign rom_data[280]=8'b00110000;
   assign rom_data[281]=8'b00101101;
   assign rom_data[282]=8'b00110000;
   assign rom_data[283]=8'b00101101;
   assign rom_data[284]=8'b00110000;
   assign rom_data[285]=8'b00101101;
   assign rom_data[286]=8'b00110000;
   assign rom_data[287]=8'b00101110;
   assign rom_data[288]=8'b00110000;
   assign rom_data[289]=8'b00101111;
   assign rom_data[290]=8'b00110000;
   assign rom_data[291]=8'b00101111;
   assign rom_data[292]=8'b00110000;
   assign rom_data[293]=8'b00110000;
   assign rom_data[294]=8'b00110000;
   assign rom_data[295]=8'b00110001;
   assign rom_data[296]=8'b00110000;
   assign rom_data[297]=8'b00110001;
   assign rom_data[298]=8'b00110000;
   assign rom_data[299]=8'b00110010;
   assign rom_data[300]=8'b00110000;
   assign rom_data[301]=8'b00110011;
   assign rom_data[302]=8'b00110000;
   assign rom_data[303]=8'b00110100;
   assign rom_data[304]=8'b00110000;
   assign rom_data[305]=8'b00110101;
   assign rom_data[306]=8'b00110000;
   assign rom_data[307]=8'b00110110;
   assign rom_data[308]=8'b00110000;
   assign rom_data[309]=8'b00110111;
   assign rom_data[310]=8'b00110000;
   assign rom_data[311]=8'b00111000;
   assign rom_data[312]=8'b00110000;
   assign rom_data[313]=8'b00111010;
   assign rom_data[314]=8'b00110000;
   assign rom_data[315]=8'b00111011;
   assign rom_data[316]=8'b00110000;
   assign rom_data[317]=8'b00111100;
   assign rom_data[318]=8'b00110000;
   assign rom_data[319]=8'b00111101;
   assign rom_data[320]=8'b00110000;
   assign rom_data[321]=8'b00111110;
   assign rom_data[322]=8'b00110000;
   assign rom_data[323]=8'b01000000;
   assign rom_data[324]=8'b00110000;
   assign rom_data[325]=8'b01000001;
   assign rom_data[326]=8'b00110000;
   assign rom_data[327]=8'b01000010;
   assign rom_data[328]=8'b00110000;
   assign rom_data[329]=8'b01000100;
   assign rom_data[330]=8'b00110000;
   assign rom_data[331]=8'b01000101;
   assign rom_data[332]=8'b00110000;
   assign rom_data[333]=8'b01000110;
   assign rom_data[334]=8'b00110001;
   assign rom_data[335]=8'b01000111;
   assign rom_data[336]=8'b00110001;
   assign rom_data[337]=8'b01001001;
   assign rom_data[338]=8'b00110001;
   assign rom_data[339]=8'b01001010;
   assign rom_data[340]=8'b00110001;
   assign rom_data[341]=8'b01001100;
   assign rom_data[342]=8'b00110001;
   assign rom_data[343]=8'b01001101;
   assign rom_data[344]=8'b00110001;
   assign rom_data[345]=8'b01001110;
   assign rom_data[346]=8'b00110001;
   assign rom_data[347]=8'b01010000;
   assign rom_data[348]=8'b00110001;
   assign rom_data[349]=8'b01010001;
   assign rom_data[350]=8'b00110001;
   assign rom_data[351]=8'b01010010;
   assign rom_data[352]=8'b00110001;
   assign rom_data[353]=8'b01010100;
   assign rom_data[354]=8'b00110001;
   assign rom_data[355]=8'b01010101;
   assign rom_data[356]=8'b00110001;
   assign rom_data[357]=8'b01010111;
   assign rom_data[358]=8'b00110001;
   assign rom_data[359]=8'b01011000;
   assign rom_data[360]=8'b00110001;
   assign rom_data[361]=8'b01011010;
   assign rom_data[362]=8'b00110001;
   assign rom_data[363]=8'b01011011;
   assign rom_data[364]=8'b00110001;
   assign rom_data[365]=8'b01011100;
   assign rom_data[366]=8'b00110001;
   assign rom_data[367]=8'b01011110;
   assign rom_data[368]=8'b00110001;
   assign rom_data[369]=8'b01011111;
   assign rom_data[370]=8'b00110001;
   assign rom_data[371]=8'b01100001;
   assign rom_data[372]=8'b00110001;
   assign rom_data[373]=8'b01100010;
   assign rom_data[374]=8'b00110001;
   assign rom_data[375]=8'b01100011;
   assign rom_data[376]=8'b00110001;
   assign rom_data[377]=8'b01100101;
   assign rom_data[378]=8'b00110001;
   assign rom_data[379]=8'b01100110;
   assign rom_data[380]=8'b00110001;
   assign rom_data[381]=8'b01100111;
   assign rom_data[382]=8'b00110001;
   assign rom_data[383]=8'b01101001;
   assign rom_data[384]=8'b00110001;
   assign rom_data[385]=8'b01101010;
   assign rom_data[386]=8'b00110001;
   assign rom_data[387]=8'b01101100;
   assign rom_data[388]=8'b00110001;
   assign rom_data[389]=8'b01101101;
   assign rom_data[390]=8'b00110001;
   assign rom_data[391]=8'b01101110;
   assign rom_data[392]=8'b00110001;
   assign rom_data[393]=8'b01110000;
   assign rom_data[394]=8'b00110001;
   assign rom_data[395]=8'b01110001;
   assign rom_data[396]=8'b00110001;
   assign rom_data[397]=8'b01110010;
   assign rom_data[398]=8'b00110001;
   assign rom_data[399]=8'b01110100;
   assign rom_data[400]=8'b00110001;
   assign rom_data[401]=8'b01110101;
   assign rom_data[402]=8'b00110001;
   assign rom_data[403]=8'b01110110;
   assign rom_data[404]=8'b00110001;
   assign rom_data[405]=8'b01110111;
   assign rom_data[406]=8'b00110001;
   assign rom_data[407]=8'b01111001;
   assign rom_data[408]=8'b00110001;
   assign rom_data[409]=8'b01111010;
   assign rom_data[410]=8'b00110001;
   assign rom_data[411]=8'b01111011;
   assign rom_data[412]=8'b00110001;
   assign rom_data[413]=8'b01111100;
   assign rom_data[414]=8'b00110001;
   assign rom_data[415]=8'b01111101;
   assign rom_data[416]=8'b00110001;
   assign rom_data[417]=8'b01111110;
   assign rom_data[418]=8'b00110010;
   assign rom_data[419]=8'b01111111;
   assign rom_data[420]=8'b00110010;
   assign rom_data[421]=8'b10000000;
   assign rom_data[422]=8'b00110010;
   assign rom_data[423]=8'b10000001;
   assign rom_data[424]=8'b00110010;
   assign rom_data[425]=8'b10000010;
   assign rom_data[426]=8'b00110010;
   assign rom_data[427]=8'b10000011;
   assign rom_data[428]=8'b00110010;
   assign rom_data[429]=8'b10000100;
   assign rom_data[430]=8'b00110010;
   assign rom_data[431]=8'b10000101;
   assign rom_data[432]=8'b00110010;
   assign rom_data[433]=8'b10000110;
   assign rom_data[434]=8'b00110010;
   assign rom_data[435]=8'b10000110;
   assign rom_data[436]=8'b00110010;
   assign rom_data[437]=8'b10000111;
   assign rom_data[438]=8'b00110010;
   assign rom_data[439]=8'b10001000;
   assign rom_data[440]=8'b00110010;
   assign rom_data[441]=8'b10001000;
   assign rom_data[442]=8'b00110010;
   assign rom_data[443]=8'b10001001;
   assign rom_data[444]=8'b00110010;
   assign rom_data[445]=8'b10001001;
   assign rom_data[446]=8'b00110010;
   assign rom_data[447]=8'b10001001;
   assign rom_data[448]=8'b00110010;
   assign rom_data[449]=8'b10001010;
   assign rom_data[450]=8'b00110010;
   assign rom_data[451]=8'b10001010;
   assign rom_data[452]=8'b00110010;
   assign rom_data[453]=8'b10001010;
   assign rom_data[454]=8'b00110010;
   assign rom_data[455]=8'b10001010;
   assign rom_data[456]=8'b00110010;
   assign rom_data[457]=8'b10001010;
   assign rom_data[458]=8'b00110010;
   assign rom_data[459]=8'b10001001;
   assign rom_data[460]=8'b00110010;
   assign rom_data[461]=8'b10001001;
   assign rom_data[462]=8'b00110010;
   assign rom_data[463]=8'b10001001;
   assign rom_data[464]=8'b00110010;
   assign rom_data[465]=8'b10001000;
   assign rom_data[466]=8'b00110010;
   assign rom_data[467]=8'b10001000;
   assign rom_data[468]=8'b00110010;
   assign rom_data[469]=8'b10000111;
   assign rom_data[470]=8'b00110010;
   assign rom_data[471]=8'b10000111;
   assign rom_data[472]=8'b00110010;
   assign rom_data[473]=8'b10000110;
   assign rom_data[474]=8'b00110010;
   assign rom_data[475]=8'b10000101;
   assign rom_data[476]=8'b00110010;
   assign rom_data[477]=8'b10000100;
   assign rom_data[478]=8'b00110010;
   assign rom_data[479]=8'b10000011;
   assign rom_data[480]=8'b00110010;
   assign rom_data[481]=8'b10000011;
   assign rom_data[482]=8'b00110011;
   assign rom_data[483]=8'b10000010;
   assign rom_data[484]=8'b00110011;
   assign rom_data[485]=8'b10000001;
   assign rom_data[486]=8'b00110011;
   assign rom_data[487]=8'b10000000;
   assign rom_data[488]=8'b00110011;
   assign rom_data[489]=8'b01111110;
   assign rom_data[490]=8'b00110011;
   assign rom_data[491]=8'b01111101;
   assign rom_data[492]=8'b00110011;
   assign rom_data[493]=8'b01111100;
   assign rom_data[494]=8'b00110011;
   assign rom_data[495]=8'b01111011;
   assign rom_data[496]=8'b00110011;
   assign rom_data[497]=8'b01111010;
   assign rom_data[498]=8'b00110011;
   assign rom_data[499]=8'b01111001;
   assign rom_data[500]=8'b00110011;
   assign rom_data[501]=8'b01110111;
   assign rom_data[502]=8'b00110011;
   assign rom_data[503]=8'b01110110;
   assign rom_data[504]=8'b00110011;
   assign rom_data[505]=8'b01110101;
   assign rom_data[506]=8'b00110011;
   assign rom_data[507]=8'b01110100;
   assign rom_data[508]=8'b00110011;
   assign rom_data[509]=8'b01110010;
   assign rom_data[510]=8'b00110011;
   assign rom_data[511]=8'b01110001;
   assign rom_data[512]=8'b00110011;
   assign rom_data[513]=8'b01110000;
   assign rom_data[514]=8'b00110011;
   assign rom_data[515]=8'b01101110;
   assign rom_data[516]=8'b00110011;
   assign rom_data[517]=8'b01101101;
   assign rom_data[518]=8'b00110011;
   assign rom_data[519]=8'b01101100;
   assign rom_data[520]=8'b00110011;
   assign rom_data[521]=8'b01101010;
   assign rom_data[522]=8'b00110011;
   assign rom_data[523]=8'b01101001;
   assign rom_data[524]=8'b00110011;
   assign rom_data[525]=8'b01101000;
   assign rom_data[526]=8'b00110011;
   assign rom_data[527]=8'b01100110;
   assign rom_data[528]=8'b00110011;
   assign rom_data[529]=8'b01100101;
   assign rom_data[530]=8'b00110011;
   assign rom_data[531]=8'b01100011;
   assign rom_data[532]=8'b00110011;
   assign rom_data[533]=8'b01100010;
   assign rom_data[534]=8'b00110011;
   assign rom_data[535]=8'b01100001;
   assign rom_data[536]=8'b00110011;
   assign rom_data[537]=8'b01011111;
   assign rom_data[538]=8'b00110011;
   assign rom_data[539]=8'b01011110;
   assign rom_data[540]=8'b00110011;
   assign rom_data[541]=8'b01011100;
   assign rom_data[542]=8'b00110011;
   assign rom_data[543]=8'b01011011;
   assign rom_data[544]=8'b00110011;
   assign rom_data[545]=8'b01011001;
   assign rom_data[546]=8'b00110011;
   assign rom_data[547]=8'b01011000;
   assign rom_data[548]=8'b00110011;
   assign rom_data[549]=8'b01010111;
   assign rom_data[550]=8'b00110011;
   assign rom_data[551]=8'b01010101;
   assign rom_data[552]=8'b00110011;
   assign rom_data[553]=8'b01010100;
   assign rom_data[554]=8'b00110011;
   assign rom_data[555]=8'b01010010;
   assign rom_data[556]=8'b00110011;
   assign rom_data[557]=8'b01010001;
   assign rom_data[558]=8'b00110011;
   assign rom_data[559]=8'b01010000;
   assign rom_data[560]=8'b00110011;
   assign rom_data[561]=8'b01001110;
   assign rom_data[562]=8'b00110011;
   assign rom_data[563]=8'b01001101;
   assign rom_data[564]=8'b00110100;
   assign rom_data[565]=8'b01001100;
   assign rom_data[566]=8'b00110100;
   assign rom_data[567]=8'b01001010;
   assign rom_data[568]=8'b00110100;
   assign rom_data[569]=8'b01001001;
   assign rom_data[570]=8'b00110100;
   assign rom_data[571]=8'b01001000;
   assign rom_data[572]=8'b00110100;
   assign rom_data[573]=8'b01000110;
   assign rom_data[574]=8'b00110100;
   assign rom_data[575]=8'b01000101;
   assign rom_data[576]=8'b00110100;
   assign rom_data[577]=8'b01000100;
   assign rom_data[578]=8'b00110100;
   assign rom_data[579]=8'b01000010;
   assign rom_data[580]=8'b00110100;
   assign rom_data[581]=8'b01000001;
   assign rom_data[582]=8'b00110100;
   assign rom_data[583]=8'b01000000;
   assign rom_data[584]=8'b00110100;
   assign rom_data[585]=8'b00111111;
   assign rom_data[586]=8'b00110100;
   assign rom_data[587]=8'b00111101;
   assign rom_data[588]=8'b00110100;
   assign rom_data[589]=8'b00111100;
   assign rom_data[590]=8'b00110100;
   assign rom_data[591]=8'b00111011;
   assign rom_data[592]=8'b00110100;
   assign rom_data[593]=8'b00111010;
   assign rom_data[594]=8'b00110100;
   assign rom_data[595]=8'b00111001;
   assign rom_data[596]=8'b00110100;
   assign rom_data[597]=8'b00111000;
   assign rom_data[598]=8'b00110100;
   assign rom_data[599]=8'b00110110;
   assign rom_data[600]=8'b00110100;
   assign rom_data[601]=8'b00110101;
   assign rom_data[602]=8'b00110100;
   assign rom_data[603]=8'b00110100;
   assign rom_data[604]=8'b00110100;
   assign rom_data[605]=8'b00110011;
   assign rom_data[606]=8'b00110100;
   assign rom_data[607]=8'b00110011;
   assign rom_data[608]=8'b00110100;
   assign rom_data[609]=8'b00110010;
   assign rom_data[610]=8'b00110100;
   assign rom_data[611]=8'b00110001;
   assign rom_data[612]=8'b00110100;
   assign rom_data[613]=8'b00110000;
   assign rom_data[614]=8'b00110100;
   assign rom_data[615]=8'b00101111;
   assign rom_data[616]=8'b00110100;
   assign rom_data[617]=8'b00101111;
   assign rom_data[618]=8'b00110100;
   assign rom_data[619]=8'b00101110;
   assign rom_data[620]=8'b00110100;
   assign rom_data[621]=8'b00101110;
   assign rom_data[622]=8'b00110100;
   assign rom_data[623]=8'b00101101;
   assign rom_data[624]=8'b00110100;
   assign rom_data[625]=8'b00101101;
   assign rom_data[626]=8'b00110100;
   assign rom_data[627]=8'b00101100;
   assign rom_data[628]=8'b00110100;
   assign rom_data[629]=8'b00101100;
   assign rom_data[630]=8'b00110100;
   assign rom_data[631]=8'b00101100;
   assign rom_data[632]=8'b00110100;
   assign rom_data[633]=8'b00101100;
   assign rom_data[634]=8'b00110100;
   assign rom_data[635]=8'b00101100;
   assign rom_data[636]=8'b00110101;
   assign rom_data[637]=8'b00101100;
   assign rom_data[638]=8'b00110101;
   assign rom_data[639]=8'b00101100;
   assign rom_data[640]=8'b00110101;
   assign rom_data[641]=8'b00101101;
   assign rom_data[642]=8'b00110101;
   assign rom_data[643]=8'b00101101;
   assign rom_data[644]=8'b00110101;
   assign rom_data[645]=8'b00101101;
   assign rom_data[646]=8'b00110101;
   assign rom_data[647]=8'b00101110;
   assign rom_data[648]=8'b00110101;
   assign rom_data[649]=8'b00101111;
   assign rom_data[650]=8'b00110101;
   assign rom_data[651]=8'b00101111;
   assign rom_data[652]=8'b00110101;
   assign rom_data[653]=8'b00110000;
   assign rom_data[654]=8'b00110101;
   assign rom_data[655]=8'b00110001;
   assign rom_data[656]=8'b00110101;
   assign rom_data[657]=8'b00110001;
   assign rom_data[658]=8'b00110101;
   assign rom_data[659]=8'b00110010;
   assign rom_data[660]=8'b00110101;
   assign rom_data[661]=8'b00110011;
   assign rom_data[662]=8'b00110101;
   assign rom_data[663]=8'b00110100;
   assign rom_data[664]=8'b00110101;
   assign rom_data[665]=8'b00110101;
   assign rom_data[666]=8'b00110101;
   assign rom_data[667]=8'b00110110;
   assign rom_data[668]=8'b00110101;
   assign rom_data[669]=8'b00110111;
   assign rom_data[670]=8'b00110101;
   assign rom_data[671]=8'b00111000;
   assign rom_data[672]=8'b00110101;
   assign rom_data[673]=8'b00111010;
   assign rom_data[674]=8'b00110101;
   assign rom_data[675]=8'b00111011;
   assign rom_data[676]=8'b00110101;
   assign rom_data[677]=8'b00111100;
   assign rom_data[678]=8'b00110101;
   assign rom_data[679]=8'b00111101;
   assign rom_data[680]=8'b00110101;
   assign rom_data[681]=8'b00111110;
   assign rom_data[682]=8'b00110101;
   assign rom_data[683]=8'b01000000;
   assign rom_data[684]=8'b00110101;
   assign rom_data[685]=8'b01000001;
   assign rom_data[686]=8'b00110101;
   assign rom_data[687]=8'b01000010;
   assign rom_data[688]=8'b00110101;
   assign rom_data[689]=8'b01000100;
   assign rom_data[690]=8'b00110101;
   assign rom_data[691]=8'b01000101;
   assign rom_data[692]=8'b00110101;
   assign rom_data[693]=8'b01000110;
   assign rom_data[694]=8'b00110101;
   assign rom_data[695]=8'b01000111;
   assign rom_data[696]=8'b00110101;
   assign rom_data[697]=8'b01001001;
   assign rom_data[698]=8'b00110101;
   assign rom_data[699]=8'b01001010;
   assign rom_data[700]=8'b00110101;
   assign rom_data[701]=8'b01001100;
   assign rom_data[702]=8'b00110101;
   assign rom_data[703]=8'b01001101;
   assign rom_data[704]=8'b00110101;
   assign rom_data[705]=8'b01001110;
   assign rom_data[706]=8'b00110101;
   assign rom_data[707]=8'b01010000;
   assign rom_data[708]=8'b00110101;
   assign rom_data[709]=8'b01010001;
   assign rom_data[710]=8'b00110110;
   assign rom_data[711]=8'b01010010;
   assign rom_data[712]=8'b00110110;
   assign rom_data[713]=8'b01010100;
   assign rom_data[714]=8'b00110110;
   assign rom_data[715]=8'b01010101;
   assign rom_data[716]=8'b00110110;
   assign rom_data[717]=8'b01010111;
   assign rom_data[718]=8'b00110110;
   assign rom_data[719]=8'b01011000;
   assign rom_data[720]=8'b00110110;
   assign rom_data[721]=8'b01011010;
   assign rom_data[722]=8'b00110110;
   assign rom_data[723]=8'b01011011;
   assign rom_data[724]=8'b00110110;
   assign rom_data[725]=8'b01011100;
   assign rom_data[726]=8'b00110110;
   assign rom_data[727]=8'b01011110;
   assign rom_data[728]=8'b00110110;
   assign rom_data[729]=8'b01011111;
   assign rom_data[730]=8'b00110110;
   assign rom_data[731]=8'b01100001;
   assign rom_data[732]=8'b00110110;
   assign rom_data[733]=8'b01100010;
   assign rom_data[734]=8'b00110110;
   assign rom_data[735]=8'b01100011;
   assign rom_data[736]=8'b00110110;
   assign rom_data[737]=8'b01100101;
   assign rom_data[738]=8'b00110110;
   assign rom_data[739]=8'b01100110;
   assign rom_data[740]=8'b00110110;
   assign rom_data[741]=8'b01100111;
   assign rom_data[742]=8'b00110110;
   assign rom_data[743]=8'b01101001;
   assign rom_data[744]=8'b00110110;
   assign rom_data[745]=8'b01101010;
   assign rom_data[746]=8'b00110110;
   assign rom_data[747]=8'b01101100;
   assign rom_data[748]=8'b00110110;
   assign rom_data[749]=8'b01101101;
   assign rom_data[750]=8'b00110110;
   assign rom_data[751]=8'b01101110;
   assign rom_data[752]=8'b00110110;
   assign rom_data[753]=8'b01110000;
   assign rom_data[754]=8'b00110110;
   assign rom_data[755]=8'b01110001;
   assign rom_data[756]=8'b00110110;
   assign rom_data[757]=8'b01110010;
   assign rom_data[758]=8'b00110110;
   assign rom_data[759]=8'b01110100;
   assign rom_data[760]=8'b00110110;
   assign rom_data[761]=8'b01110101;
   assign rom_data[762]=8'b00110110;
   assign rom_data[763]=8'b01110110;
   assign rom_data[764]=8'b00110110;
   assign rom_data[765]=8'b01110111;
   assign rom_data[766]=8'b00110110;
   assign rom_data[767]=8'b01111001;
   assign rom_data[768]=8'b00110110;
   assign rom_data[769]=8'b01111010;
   assign rom_data[770]=8'b00110110;
   assign rom_data[771]=8'b01111011;
   assign rom_data[772]=8'b00110110;
   assign rom_data[773]=8'b01111100;
   assign rom_data[774]=8'b00110110;
   assign rom_data[775]=8'b01111101;
   assign rom_data[776]=8'b00110110;
   assign rom_data[777]=8'b01111110;
   assign rom_data[778]=8'b00110110;
   assign rom_data[779]=8'b01111111;
   assign rom_data[780]=8'b00110110;
   assign rom_data[781]=8'b10000000;
   assign rom_data[782]=8'b00110110;
   assign rom_data[783]=8'b10000001;
   assign rom_data[784]=8'b00110110;
   assign rom_data[785]=8'b10000010;
   assign rom_data[786]=8'b00110110;
   assign rom_data[787]=8'b10000011;
   assign rom_data[788]=8'b00110110;
   assign rom_data[789]=8'b10000100;
   assign rom_data[790]=8'b00110111;
   assign rom_data[791]=8'b10000101;
   assign rom_data[792]=8'b00110111;
   assign rom_data[793]=8'b10000110;
   assign rom_data[794]=8'b00110111;
   assign rom_data[795]=8'b10000110;
   assign rom_data[796]=8'b00110111;
   assign rom_data[797]=8'b10000111;
   assign rom_data[798]=8'b00110111;
   assign rom_data[799]=8'b10001000;
   assign rom_data[800]=8'b00110111;
   assign rom_data[801]=8'b10001000;
   assign rom_data[802]=8'b00110111;
   assign rom_data[803]=8'b10001001;
   assign rom_data[804]=8'b00110111;
   assign rom_data[805]=8'b10001001;
   assign rom_data[806]=8'b00110111;
   assign rom_data[807]=8'b10001001;
   assign rom_data[808]=8'b00110111;
   assign rom_data[809]=8'b10001010;
   assign rom_data[810]=8'b00110111;
   assign rom_data[811]=8'b10001010;
   assign rom_data[812]=8'b00110111;
   assign rom_data[813]=8'b10001010;
   assign rom_data[814]=8'b00110111;
   assign rom_data[815]=8'b10001010;
   assign rom_data[816]=8'b00110111;
   assign rom_data[817]=8'b10001010;
   assign rom_data[818]=8'b00110111;
   assign rom_data[819]=8'b10001001;
   assign rom_data[820]=8'b00110111;
   assign rom_data[821]=8'b10001001;
   assign rom_data[822]=8'b00110111;
   assign rom_data[823]=8'b10001001;
   assign rom_data[824]=8'b00110111;
   assign rom_data[825]=8'b10001000;
   assign rom_data[826]=8'b00110111;
   assign rom_data[827]=8'b10001000;
   assign rom_data[828]=8'b00110111;
   assign rom_data[829]=8'b10000111;
   assign rom_data[830]=8'b00110111;
   assign rom_data[831]=8'b10000111;
   assign rom_data[832]=8'b00110111;
   assign rom_data[833]=8'b10000110;
   assign rom_data[834]=8'b00110111;
   assign rom_data[835]=8'b10000101;
   assign rom_data[836]=8'b00110111;
   assign rom_data[837]=8'b10000100;
   assign rom_data[838]=8'b00110111;
   assign rom_data[839]=8'b10000011;
   assign rom_data[840]=8'b00110111;
   assign rom_data[841]=8'b10000011;
   assign rom_data[842]=8'b00110111;
   assign rom_data[843]=8'b10000010;
   assign rom_data[844]=8'b00110111;
   assign rom_data[845]=8'b10000001;
   assign rom_data[846]=8'b00110111;
   assign rom_data[847]=8'b10000000;
   assign rom_data[848]=8'b00110111;
   assign rom_data[849]=8'b01111110;
   assign rom_data[850]=8'b00110111;
   assign rom_data[851]=8'b01111101;
   assign rom_data[852]=8'b00110111;
   assign rom_data[853]=8'b01111100;
   assign rom_data[854]=8'b00110111;
   assign rom_data[855]=8'b01111011;
   assign rom_data[856]=8'b00111000;
   assign rom_data[857]=8'b01111010;
   assign rom_data[858]=8'b00111000;
   assign rom_data[859]=8'b01111001;
   assign rom_data[860]=8'b00111000;
   assign rom_data[861]=8'b01110111;
   assign rom_data[862]=8'b00111000;
   assign rom_data[863]=8'b01110110;
   assign rom_data[864]=8'b00111000;
   assign rom_data[865]=8'b01110101;
   assign rom_data[866]=8'b00111000;
   assign rom_data[867]=8'b01110100;
   assign rom_data[868]=8'b00111000;
   assign rom_data[869]=8'b01110010;
   assign rom_data[870]=8'b00111000;
   assign rom_data[871]=8'b01110001;
   assign rom_data[872]=8'b00111000;
   assign rom_data[873]=8'b01110000;
   assign rom_data[874]=8'b00111000;
   assign rom_data[875]=8'b01101110;
   assign rom_data[876]=8'b00111000;
   assign rom_data[877]=8'b01101101;
   assign rom_data[878]=8'b00111000;
   assign rom_data[879]=8'b01101100;
   assign rom_data[880]=8'b00111000;
   assign rom_data[881]=8'b01101010;
   assign rom_data[882]=8'b00111000;
   assign rom_data[883]=8'b01101001;
   assign rom_data[884]=8'b00111000;
   assign rom_data[885]=8'b01101000;
   assign rom_data[886]=8'b00111000;
   assign rom_data[887]=8'b01100110;
   assign rom_data[888]=8'b00111000;
   assign rom_data[889]=8'b01100101;
   assign rom_data[890]=8'b00111000;
   assign rom_data[891]=8'b01100011;
   assign rom_data[892]=8'b00111000;
   assign rom_data[893]=8'b01100010;
   assign rom_data[894]=8'b00111000;
   assign rom_data[895]=8'b01100001;
   assign rom_data[896]=8'b00111000;
   assign rom_data[897]=8'b01011111;
   assign rom_data[898]=8'b00111000;
   assign rom_data[899]=8'b01011110;
   assign rom_data[900]=8'b00111000;
   assign rom_data[901]=8'b01011100;
   assign rom_data[902]=8'b00111000;
   assign rom_data[903]=8'b01011011;
   assign rom_data[904]=8'b00111000;
   assign rom_data[905]=8'b01011001;
   assign rom_data[906]=8'b00111000;
   assign rom_data[907]=8'b01011000;
   assign rom_data[908]=8'b00111000;
   assign rom_data[909]=8'b01010111;
   assign rom_data[910]=8'b00111000;
   assign rom_data[911]=8'b01010101;
   assign rom_data[912]=8'b00111000;
   assign rom_data[913]=8'b01010100;
   assign rom_data[914]=8'b00111000;
   assign rom_data[915]=8'b01010010;
   assign rom_data[916]=8'b00111000;
   assign rom_data[917]=8'b01010001;
   assign rom_data[918]=8'b00111000;
   assign rom_data[919]=8'b01010000;
   assign rom_data[920]=8'b00111000;
   assign rom_data[921]=8'b01001110;
   assign rom_data[922]=8'b00111000;
   assign rom_data[923]=8'b01001101;
   assign rom_data[924]=8'b00111000;
   assign rom_data[925]=8'b01001100;
   assign rom_data[926]=8'b00111000;
   assign rom_data[927]=8'b01001010;
   assign rom_data[928]=8'b00111000;
   assign rom_data[929]=8'b01001001;
   assign rom_data[930]=8'b00111000;
   assign rom_data[931]=8'b01001000;
   assign rom_data[932]=8'b00111000;
   assign rom_data[933]=8'b01000110;
   assign rom_data[934]=8'b00111000;
   assign rom_data[935]=8'b01000101;
   assign rom_data[936]=8'b00111000;
   assign rom_data[937]=8'b01000100;
   assign rom_data[938]=8'b00111000;
   assign rom_data[939]=8'b01000010;
   assign rom_data[940]=8'b00111001;
   assign rom_data[941]=8'b01000001;
   assign rom_data[942]=8'b00111001;
   assign rom_data[943]=8'b01000000;
   assign rom_data[944]=8'b00111001;
   assign rom_data[945]=8'b00111111;
   assign rom_data[946]=8'b00111001;
   assign rom_data[947]=8'b00111101;
   assign rom_data[948]=8'b00111001;
   assign rom_data[949]=8'b00111100;
   assign rom_data[950]=8'b00111001;
   assign rom_data[951]=8'b00111011;
   assign rom_data[952]=8'b00111001;
   assign rom_data[953]=8'b00111010;
   assign rom_data[954]=8'b00111001;
   assign rom_data[955]=8'b00111001;
   assign rom_data[956]=8'b00111001;
   assign rom_data[957]=8'b00111000;
   assign rom_data[958]=8'b00111001;
   assign rom_data[959]=8'b00110110;
   assign rom_data[960]=8'b00111001;
   assign rom_data[961]=8'b00110101;
   assign rom_data[962]=8'b00111001;
   assign rom_data[963]=8'b00110100;
   assign rom_data[964]=8'b00111001;
   assign rom_data[965]=8'b00110011;
   assign rom_data[966]=8'b00111001;
   assign rom_data[967]=8'b00110011;
   assign rom_data[968]=8'b00111001;
   assign rom_data[969]=8'b00110010;
   assign rom_data[970]=8'b00111001;
   assign rom_data[971]=8'b00110001;
   assign rom_data[972]=8'b00111001;
   assign rom_data[973]=8'b00110000;
   assign rom_data[974]=8'b00111001;
   assign rom_data[975]=8'b00101111;
   assign rom_data[976]=8'b00111001;
   assign rom_data[977]=8'b00101111;
   assign rom_data[978]=8'b00111001;
   assign rom_data[979]=8'b00101110;
   assign rom_data[980]=8'b00111001;
   assign rom_data[981]=8'b00101110;
   assign rom_data[982]=8'b00111001;
   assign rom_data[983]=8'b00101101;
   assign rom_data[984]=8'b00111001;
   assign rom_data[985]=8'b00101101;
   assign rom_data[986]=8'b00111001;
   assign rom_data[987]=8'b00101100;
   assign rom_data[988]=8'b00111001;
   assign rom_data[989]=8'b00101100;
   assign rom_data[990]=8'b00111001;
   assign rom_data[991]=8'b00101100;
   assign rom_data[992]=8'b00111001;
   assign rom_data[993]=8'b00101100;
   assign rom_data[994]=8'b00111001;
   assign rom_data[995]=8'b00101100;
   assign rom_data[996]=8'b00111001;
   assign rom_data[997]=8'b00101100;
   assign rom_data[998]=8'b00111001;
   assign rom_data[999]=8'b00101100;
   assign rom_data[1000]=8'b00111001;
   assign rom_data[1001]=8'b00101101;
   assign rom_data[1002]=8'b00111001;
   assign rom_data[1003]=8'b00101101;
   assign rom_data[1004]=8'b00111001;
   assign rom_data[1005]=8'b00101101;
   assign rom_data[1006]=8'b00111001;
   assign rom_data[1007]=8'b00101110;
   assign rom_data[1008]=8'b00111010;
   assign rom_data[1009]=8'b00101111;
   assign rom_data[1010]=8'b00111010;
   assign rom_data[1011]=8'b00101111;
   assign rom_data[1012]=8'b00111010;
   assign rom_data[1013]=8'b00110000;
   assign rom_data[1014]=8'b00111010;
   assign rom_data[1015]=8'b00110001;
   assign rom_data[1016]=8'b00111010;
   assign rom_data[1017]=8'b00110001;
   assign rom_data[1018]=8'b00111010;
   assign rom_data[1019]=8'b00110010;
   assign rom_data[1020]=8'b00111010;
   assign rom_data[1021]=8'b00110011;
   assign rom_data[1022]=8'b00111010;
   assign rom_data[1023]=8'b00110100;
   assign rom_data[1024]=8'b00111010;
   assign rom_data[1025]=8'b00110101;
   assign rom_data[1026]=8'b00111010;
   assign rom_data[1027]=8'b00110110;
   assign rom_data[1028]=8'b00111010;
   assign rom_data[1029]=8'b00110111;
   assign rom_data[1030]=8'b00111010;
   assign rom_data[1031]=8'b00111000;
   assign rom_data[1032]=8'b00111010;
   assign rom_data[1033]=8'b00111010;
   assign rom_data[1034]=8'b00111010;
   assign rom_data[1035]=8'b00111011;
   assign rom_data[1036]=8'b00111010;
   assign rom_data[1037]=8'b00111100;
   assign rom_data[1038]=8'b00111010;
   assign rom_data[1039]=8'b00111101;
   assign rom_data[1040]=8'b00111010;
   assign rom_data[1041]=8'b00111110;
   assign rom_data[1042]=8'b00111010;
   assign rom_data[1043]=8'b01000000;
   assign rom_data[1044]=8'b00111010;
   assign rom_data[1045]=8'b01000001;
   assign rom_data[1046]=8'b00111010;
   assign rom_data[1047]=8'b01000010;
   assign rom_data[1048]=8'b00111010;
   assign rom_data[1049]=8'b01000100;
   assign rom_data[1050]=8'b00111010;
   assign rom_data[1051]=8'b01000101;
   assign rom_data[1052]=8'b00111010;
   assign rom_data[1053]=8'b01000110;
   assign rom_data[1054]=8'b00111010;
   assign rom_data[1055]=8'b01000111;
   assign rom_data[1056]=8'b00111010;
   assign rom_data[1057]=8'b01001001;
   assign rom_data[1058]=8'b00111010;
   assign rom_data[1059]=8'b01001010;
   assign rom_data[1060]=8'b00111010;
   assign rom_data[1061]=8'b01001100;
   assign rom_data[1062]=8'b00111010;
   assign rom_data[1063]=8'b01001101;
   assign rom_data[1064]=8'b00111010;
   assign rom_data[1065]=8'b01001110;
   assign rom_data[1066]=8'b00111010;
   assign rom_data[1067]=8'b01010000;
   assign rom_data[1068]=8'b00111010;
   assign rom_data[1069]=8'b01010001;
   assign rom_data[1070]=8'b00111010;
   assign rom_data[1071]=8'b01010010;
   assign rom_data[1072]=8'b00111010;
   assign rom_data[1073]=8'b01010100;
   assign rom_data[1074]=8'b00111010;
   assign rom_data[1075]=8'b01010101;
   assign rom_data[1076]=8'b00111010;
   assign rom_data[1077]=8'b01010111;
   assign rom_data[1078]=8'b00111010;
   assign rom_data[1079]=8'b01011000;
   assign rom_data[1080]=8'b00111010;
   assign rom_data[1081]=8'b01011010;
   assign rom_data[1082]=8'b00111010;
   assign rom_data[1083]=8'b01011011;
   assign rom_data[1084]=8'b00111010;
   assign rom_data[1085]=8'b01011100;
   assign rom_data[1086]=8'b00111011;
   assign rom_data[1087]=8'b01011110;
   assign rom_data[1088]=8'b00111011;
   assign rom_data[1089]=8'b01011111;
   assign rom_data[1090]=8'b00111011;
   assign rom_data[1091]=8'b01100001;
   assign rom_data[1092]=8'b00111011;
   assign rom_data[1093]=8'b01100010;
   assign rom_data[1094]=8'b00111011;
   assign rom_data[1095]=8'b01100011;
   assign rom_data[1096]=8'b00111011;
   assign rom_data[1097]=8'b01100101;
   assign rom_data[1098]=8'b00111011;
   assign rom_data[1099]=8'b01100110;
   assign rom_data[1100]=8'b00111011;
   assign rom_data[1101]=8'b01100111;
   assign rom_data[1102]=8'b00111011;
   assign rom_data[1103]=8'b01101001;
   assign rom_data[1104]=8'b00111011;
   assign rom_data[1105]=8'b01101010;
   assign rom_data[1106]=8'b00111011;
   assign rom_data[1107]=8'b01101100;
   assign rom_data[1108]=8'b00111011;
   assign rom_data[1109]=8'b01101101;
   assign rom_data[1110]=8'b00111011;
   assign rom_data[1111]=8'b01101110;
   assign rom_data[1112]=8'b00111011;
   assign rom_data[1113]=8'b01110000;
   assign rom_data[1114]=8'b00111011;
   assign rom_data[1115]=8'b01110001;
   assign rom_data[1116]=8'b00111011;
   assign rom_data[1117]=8'b01110010;
   assign rom_data[1118]=8'b00111011;
   assign rom_data[1119]=8'b01110100;
   assign rom_data[1120]=8'b00111011;
   assign rom_data[1121]=8'b01110101;
   assign rom_data[1122]=8'b00111011;
   assign rom_data[1123]=8'b01110110;
   assign rom_data[1124]=8'b00111011;
   assign rom_data[1125]=8'b01110111;
   assign rom_data[1126]=8'b00111011;
   assign rom_data[1127]=8'b01111001;
   assign rom_data[1128]=8'b00111011;
   assign rom_data[1129]=8'b01111010;
   assign rom_data[1130]=8'b00111011;
   assign rom_data[1131]=8'b01111011;
   assign rom_data[1132]=8'b00111011;
   assign rom_data[1133]=8'b01111100;
   assign rom_data[1134]=8'b00111011;
   assign rom_data[1135]=8'b01111101;
   assign rom_data[1136]=8'b00111011;
   assign rom_data[1137]=8'b01111110;
   assign rom_data[1138]=8'b00111011;
   assign rom_data[1139]=8'b01111111;
   assign rom_data[1140]=8'b00111011;
   assign rom_data[1141]=8'b10000000;
   assign rom_data[1142]=8'b00111011;
   assign rom_data[1143]=8'b10000001;
   assign rom_data[1144]=8'b00111011;
   assign rom_data[1145]=8'b10000010;
   assign rom_data[1146]=8'b00111011;
   assign rom_data[1147]=8'b10000011;
   assign rom_data[1148]=8'b00111011;
   assign rom_data[1149]=8'b10000100;
   assign rom_data[1150]=8'b00111011;
   assign rom_data[1151]=8'b10000101;
   assign rom_data[1152]=8'b00111011;
   assign rom_data[1153]=8'b10000110;
   assign rom_data[1154]=8'b00111011;
   assign rom_data[1155]=8'b10000110;
   assign rom_data[1156]=8'b00111011;
   assign rom_data[1157]=8'b10000111;
   assign rom_data[1158]=8'b00111011;
   assign rom_data[1159]=8'b10001000;
   assign rom_data[1160]=8'b00111011;
   assign rom_data[1161]=8'b10001000;
   assign rom_data[1162]=8'b00111011;
   assign rom_data[1163]=8'b10001001;
   assign rom_data[1164]=8'b00111100;
   assign rom_data[1165]=8'b10001001;
   assign rom_data[1166]=8'b00111100;
   assign rom_data[1167]=8'b10001001;
   assign rom_data[1168]=8'b00111100;
   assign rom_data[1169]=8'b10001010;
   assign rom_data[1170]=8'b00111100;
   assign rom_data[1171]=8'b10001010;
   assign rom_data[1172]=8'b00111100;
   assign rom_data[1173]=8'b10001010;
   assign rom_data[1174]=8'b00111100;
   assign rom_data[1175]=8'b10001010;
   assign rom_data[1176]=8'b00111100;
   assign rom_data[1177]=8'b10001010;
   assign rom_data[1178]=8'b00111100;
   assign rom_data[1179]=8'b10001001;
   assign rom_data[1180]=8'b00111100;
   assign rom_data[1181]=8'b10001001;
   assign rom_data[1182]=8'b00111100;
   assign rom_data[1183]=8'b10001001;
   assign rom_data[1184]=8'b00111100;
   assign rom_data[1185]=8'b10001000;
   assign rom_data[1186]=8'b00111100;
   assign rom_data[1187]=8'b10001000;
   assign rom_data[1188]=8'b00111100;
   assign rom_data[1189]=8'b10000111;
   assign rom_data[1190]=8'b00111100;
   assign rom_data[1191]=8'b10000111;
   assign rom_data[1192]=8'b00111100;
   assign rom_data[1193]=8'b10000110;
   assign rom_data[1194]=8'b00111100;
   assign rom_data[1195]=8'b10000101;
   assign rom_data[1196]=8'b00111100;
   assign rom_data[1197]=8'b10000100;
   assign rom_data[1198]=8'b00111100;
   assign rom_data[1199]=8'b10000011;
   assign rom_data[1200]=8'b00111100;
   assign rom_data[1201]=8'b10000011;
   assign rom_data[1202]=8'b00111100;
   assign rom_data[1203]=8'b10000010;
   assign rom_data[1204]=8'b00111100;
   assign rom_data[1205]=8'b10000001;
   assign rom_data[1206]=8'b00111100;
   assign rom_data[1207]=8'b10000000;
   assign rom_data[1208]=8'b00111100;
   assign rom_data[1209]=8'b01111110;
   assign rom_data[1210]=8'b00111100;
   assign rom_data[1211]=8'b01111101;
   assign rom_data[1212]=8'b00111100;
   assign rom_data[1213]=8'b01111100;
   assign rom_data[1214]=8'b00111100;
   assign rom_data[1215]=8'b01111011;
   assign rom_data[1216]=8'b00111100;
   assign rom_data[1217]=8'b01111010;
   assign rom_data[1218]=8'b00111100;
   assign rom_data[1219]=8'b01111001;
   assign rom_data[1220]=8'b00111100;
   assign rom_data[1221]=8'b01110111;
   assign rom_data[1222]=8'b00111100;
   assign rom_data[1223]=8'b01110110;
   assign rom_data[1224]=8'b00111100;
   assign rom_data[1225]=8'b01110101;
   assign rom_data[1226]=8'b00111100;
   assign rom_data[1227]=8'b01110100;
   assign rom_data[1228]=8'b00111100;
   assign rom_data[1229]=8'b01110010;
   assign rom_data[1230]=8'b00111100;
   assign rom_data[1231]=8'b01110001;
   assign rom_data[1232]=8'b00111101;
   assign rom_data[1233]=8'b01110000;
   assign rom_data[1234]=8'b00111101;
   assign rom_data[1235]=8'b01101110;
   assign rom_data[1236]=8'b00111101;
   assign rom_data[1237]=8'b01101101;
   assign rom_data[1238]=8'b00111101;
   assign rom_data[1239]=8'b01101100;
   assign rom_data[1240]=8'b00111101;
   assign rom_data[1241]=8'b01101010;
   assign rom_data[1242]=8'b00111101;
   assign rom_data[1243]=8'b01101001;
   assign rom_data[1244]=8'b00111101;
   assign rom_data[1245]=8'b01100111;
   assign rom_data[1246]=8'b00111101;
   assign rom_data[1247]=8'b01100110;
   assign rom_data[1248]=8'b00111101;
   assign rom_data[1249]=8'b01100101;
   assign rom_data[1250]=8'b00111101;
   assign rom_data[1251]=8'b01100011;
   assign rom_data[1252]=8'b00111101;
   assign rom_data[1253]=8'b01100010;
   assign rom_data[1254]=8'b00111101;
   assign rom_data[1255]=8'b01100001;
   assign rom_data[1256]=8'b00111101;
   assign rom_data[1257]=8'b01011111;
   assign rom_data[1258]=8'b00111101;
   assign rom_data[1259]=8'b01011110;
   assign rom_data[1260]=8'b00111101;
   assign rom_data[1261]=8'b01011100;
   assign rom_data[1262]=8'b00111101;
   assign rom_data[1263]=8'b01011011;
   assign rom_data[1264]=8'b00111101;
   assign rom_data[1265]=8'b01011001;
   assign rom_data[1266]=8'b00111101;
   assign rom_data[1267]=8'b01011000;
   assign rom_data[1268]=8'b00111101;
   assign rom_data[1269]=8'b01010111;
   assign rom_data[1270]=8'b00111101;
   assign rom_data[1271]=8'b01010101;
   assign rom_data[1272]=8'b00111101;
   assign rom_data[1273]=8'b01010100;
   assign rom_data[1274]=8'b00111101;
   assign rom_data[1275]=8'b01010010;
   assign rom_data[1276]=8'b00111101;
   assign rom_data[1277]=8'b01010001;
   assign rom_data[1278]=8'b00111101;
   assign rom_data[1279]=8'b01010000;
   assign rom_data[1280]=8'b00111101;
   assign rom_data[1281]=8'b01001110;
   assign rom_data[1282]=8'b00111101;
   assign rom_data[1283]=8'b01001101;
   assign rom_data[1284]=8'b00111101;
   assign rom_data[1285]=8'b01001100;
   assign rom_data[1286]=8'b00111101;
   assign rom_data[1287]=8'b01001010;
   assign rom_data[1288]=8'b00111101;
   assign rom_data[1289]=8'b01001001;
   assign rom_data[1290]=8'b00111101;
   assign rom_data[1291]=8'b01001000;
   assign rom_data[1292]=8'b00111101;
   assign rom_data[1293]=8'b01000110;
   assign rom_data[1294]=8'b00111101;
   assign rom_data[1295]=8'b01000101;
   assign rom_data[1296]=8'b00111101;
   assign rom_data[1297]=8'b01000100;
   assign rom_data[1298]=8'b00111101;
   assign rom_data[1299]=8'b01000010;
   assign rom_data[1300]=8'b00111101;
   assign rom_data[1301]=8'b01000001;
   assign rom_data[1302]=8'b00111101;
   assign rom_data[1303]=8'b01000000;
   assign rom_data[1304]=8'b00111101;
   assign rom_data[1305]=8'b00111111;
   assign rom_data[1306]=8'b00111101;
   assign rom_data[1307]=8'b00111101;
   assign rom_data[1308]=8'b00111101;
   assign rom_data[1309]=8'b00111100;
   assign rom_data[1310]=8'b00111101;
   assign rom_data[1311]=8'b00111011;
   assign rom_data[1312]=8'b00111101;
   assign rom_data[1313]=8'b00111010;
   assign rom_data[1314]=8'b00111101;
   assign rom_data[1315]=8'b00111001;
   assign rom_data[1316]=8'b00111110;
   assign rom_data[1317]=8'b00111000;
   assign rom_data[1318]=8'b00111110;
   assign rom_data[1319]=8'b00110110;
   assign rom_data[1320]=8'b00111110;
   assign rom_data[1321]=8'b00110101;
   assign rom_data[1322]=8'b00111110;
   assign rom_data[1323]=8'b00110100;
   assign rom_data[1324]=8'b00111110;
   assign rom_data[1325]=8'b00110011;
   assign rom_data[1326]=8'b00111110;
   assign rom_data[1327]=8'b00110011;
   assign rom_data[1328]=8'b00111110;
   assign rom_data[1329]=8'b00110010;
   assign rom_data[1330]=8'b00111110;
   assign rom_data[1331]=8'b00110001;
   assign rom_data[1332]=8'b00111110;
   assign rom_data[1333]=8'b00110000;
   assign rom_data[1334]=8'b00111110;
   assign rom_data[1335]=8'b00101111;
   assign rom_data[1336]=8'b00111110;
   assign rom_data[1337]=8'b00101111;
   assign rom_data[1338]=8'b00111110;
   assign rom_data[1339]=8'b00101110;
   assign rom_data[1340]=8'b00111110;
   assign rom_data[1341]=8'b00101110;
   assign rom_data[1342]=8'b00111110;
   assign rom_data[1343]=8'b00101101;
   assign rom_data[1344]=8'b00111110;
   assign rom_data[1345]=8'b00101101;
   assign rom_data[1346]=8'b00111110;
   assign rom_data[1347]=8'b00101100;
   assign rom_data[1348]=8'b00111110;
   assign rom_data[1349]=8'b00101100;
   assign rom_data[1350]=8'b00111110;
   assign rom_data[1351]=8'b00101100;
   assign rom_data[1352]=8'b00111110;
   assign rom_data[1353]=8'b00101100;
   assign rom_data[1354]=8'b00111110;
   assign rom_data[1355]=8'b00101100;
   assign rom_data[1356]=8'b00111110;
   assign rom_data[1357]=8'b00101100;
   assign rom_data[1358]=8'b00111110;
   assign rom_data[1359]=8'b00101100;
   assign rom_data[1360]=8'b00111110;
   assign rom_data[1361]=8'b00101101;
   assign rom_data[1362]=8'b00111110;
   assign rom_data[1363]=8'b00101101;
   assign rom_data[1364]=8'b00111110;
   assign rom_data[1365]=8'b00101101;
   assign rom_data[1366]=8'b00111110;
   assign rom_data[1367]=8'b00101110;
   assign rom_data[1368]=8'b00111110;
   assign rom_data[1369]=8'b00101111;
   assign rom_data[1370]=8'b00111110;
   assign rom_data[1371]=8'b00101111;
   assign rom_data[1372]=8'b00111110;
   assign rom_data[1373]=8'b00110000;
   assign rom_data[1374]=8'b00111110;
   assign rom_data[1375]=8'b00110001;
   assign rom_data[1376]=8'b00111110;
   assign rom_data[1377]=8'b00110001;
   assign rom_data[1378]=8'b00111110;
   assign rom_data[1379]=8'b00110010;
   assign rom_data[1380]=8'b00111110;
   assign rom_data[1381]=8'b00110011;
   assign rom_data[1382]=8'b00111111;
   assign rom_data[1383]=8'b00110100;
   assign rom_data[1384]=8'b00111111;
   assign rom_data[1385]=8'b00110101;
   assign rom_data[1386]=8'b00111111;
   assign rom_data[1387]=8'b00110110;
   assign rom_data[1388]=8'b00111111;
   assign rom_data[1389]=8'b00110111;
   assign rom_data[1390]=8'b00111111;
   assign rom_data[1391]=8'b00111000;
   assign rom_data[1392]=8'b00111111;
   assign rom_data[1393]=8'b00111010;
   assign rom_data[1394]=8'b00111111;
   assign rom_data[1395]=8'b00111011;
   assign rom_data[1396]=8'b00111111;
   assign rom_data[1397]=8'b00111100;
   assign rom_data[1398]=8'b00111111;
   assign rom_data[1399]=8'b00111101;
   assign rom_data[1400]=8'b00111111;
   assign rom_data[1401]=8'b00111110;
   assign rom_data[1402]=8'b00111111;
   assign rom_data[1403]=8'b01000000;
   assign rom_data[1404]=8'b00111111;
   assign rom_data[1405]=8'b01000001;
   assign rom_data[1406]=8'b00111111;
   assign rom_data[1407]=8'b01000010;
   assign rom_data[1408]=8'b00111111;
   assign rom_data[1409]=8'b01000100;
   assign rom_data[1410]=8'b00111111;
   assign rom_data[1411]=8'b01000101;
   assign rom_data[1412]=8'b00111111;
   assign rom_data[1413]=8'b01000110;
   assign rom_data[1414]=8'b00111111;
   assign rom_data[1415]=8'b01000111;
   assign rom_data[1416]=8'b00111111;
   assign rom_data[1417]=8'b01001001;
   assign rom_data[1418]=8'b00111111;
   assign rom_data[1419]=8'b01001010;
   assign rom_data[1420]=8'b00111111;
   assign rom_data[1421]=8'b01001100;
   assign rom_data[1422]=8'b00111111;
   assign rom_data[1423]=8'b01001101;
   assign rom_data[1424]=8'b00111111;
   assign rom_data[1425]=8'b01001110;
   assign rom_data[1426]=8'b00111111;
   assign rom_data[1427]=8'b01010000;
   assign rom_data[1428]=8'b00111111;
   assign rom_data[1429]=8'b01010001;
   assign rom_data[1430]=8'b00111111;
   assign rom_data[1431]=8'b01010010;
   assign rom_data[1432]=8'b00111111;
   assign rom_data[1433]=8'b01010100;
   assign rom_data[1434]=8'b00111111;
   assign rom_data[1435]=8'b01010101;
   assign rom_data[1436]=8'b00111111;
   assign rom_data[1437]=8'b01010111;
   assign rom_data[1438]=8'b00111111;
   assign rom_data[1439]=8'b01011000;
   assign rom_data[1440]=8'b00111111;
   assign rom_data[1441]=8'b01011010;
   assign rom_data[1442]=8'b00111111;
   assign rom_data[1443]=8'b01011011;
   assign rom_data[1444]=8'b00111111;
   assign rom_data[1445]=8'b01011100;
   assign rom_data[1446]=8'b00111111;
   assign rom_data[1447]=8'b01011110;
   assign rom_data[1448]=8'b00111111;
   assign rom_data[1449]=8'b01011111;
   assign rom_data[1450]=8'b00111111;
   assign rom_data[1451]=8'b01100001;
   assign rom_data[1452]=8'b00111111;
   assign rom_data[1453]=8'b01100010;
   assign rom_data[1454]=8'b00111111;
   assign rom_data[1455]=8'b01100011;
   assign rom_data[1456]=8'b00111111;
   assign rom_data[1457]=8'b01100101;
   assign rom_data[1458]=8'b00111111;
   assign rom_data[1459]=8'b01100110;
   assign rom_data[1460]=8'b00111111;
   assign rom_data[1461]=8'b01100111;
   assign rom_data[1462]=8'b00111111;
   assign rom_data[1463]=8'b01101001;
   assign rom_data[1464]=8'b01000000;
   assign rom_data[1465]=8'b01101010;
   assign rom_data[1466]=8'b01000000;
   assign rom_data[1467]=8'b01101100;
   assign rom_data[1468]=8'b01000000;
   assign rom_data[1469]=8'b01101101;
   assign rom_data[1470]=8'b01000000;
   assign rom_data[1471]=8'b01101110;
   assign rom_data[1472]=8'b01000000;
   assign rom_data[1473]=8'b01110000;
   assign rom_data[1474]=8'b01000000;
   assign rom_data[1475]=8'b01110001;
   assign rom_data[1476]=8'b01000000;
   assign rom_data[1477]=8'b01110010;
   assign rom_data[1478]=8'b01000000;
   assign rom_data[1479]=8'b01110100;
   assign rom_data[1480]=8'b01000000;
   assign rom_data[1481]=8'b01110101;
   assign rom_data[1482]=8'b01000000;
   assign rom_data[1483]=8'b01110110;
   assign rom_data[1484]=8'b01000000;
   assign rom_data[1485]=8'b01110111;
   assign rom_data[1486]=8'b01000000;
   assign rom_data[1487]=8'b01111001;
   assign rom_data[1488]=8'b01000000;
   assign rom_data[1489]=8'b01111010;
   assign rom_data[1490]=8'b01000000;
   assign rom_data[1491]=8'b01111011;
   assign rom_data[1492]=8'b01000000;
   assign rom_data[1493]=8'b01111100;
   assign rom_data[1494]=8'b01000000;
   assign rom_data[1495]=8'b01111101;
   assign rom_data[1496]=8'b01000000;
   assign rom_data[1497]=8'b01111110;
   assign rom_data[1498]=8'b01000000;
   assign rom_data[1499]=8'b01111111;
   assign rom_data[1500]=8'b01000000;
   assign rom_data[1501]=8'b10000000;
   assign rom_data[1502]=8'b01000000;
   assign rom_data[1503]=8'b10000001;
   assign rom_data[1504]=8'b01000000;
   assign rom_data[1505]=8'b10000010;
   assign rom_data[1506]=8'b01000000;
   assign rom_data[1507]=8'b10000011;
   assign rom_data[1508]=8'b01000000;
   assign rom_data[1509]=8'b10000100;
   assign rom_data[1510]=8'b01000000;
   assign rom_data[1511]=8'b10000101;
   assign rom_data[1512]=8'b01000000;
   assign rom_data[1513]=8'b10000110;
   assign rom_data[1514]=8'b01000000;
   assign rom_data[1515]=8'b10000110;
   assign rom_data[1516]=8'b01000000;
   assign rom_data[1517]=8'b10000111;
   assign rom_data[1518]=8'b01000000;
   assign rom_data[1519]=8'b10001000;
   assign rom_data[1520]=8'b01000000;
   assign rom_data[1521]=8'b10001000;
   assign rom_data[1522]=8'b01000000;
   assign rom_data[1523]=8'b10001001;
   assign rom_data[1524]=8'b01000000;
   assign rom_data[1525]=8'b10001001;
   assign rom_data[1526]=8'b01000000;
   assign rom_data[1527]=8'b10001001;
   assign rom_data[1528]=8'b01000000;
   assign rom_data[1529]=8'b10001010;
   assign rom_data[1530]=8'b01000000;
   assign rom_data[1531]=8'b10001010;
   assign rom_data[1532]=8'b01000000;
   assign rom_data[1533]=8'b10001010;
   assign rom_data[1534]=8'b01000000;
   assign rom_data[1535]=8'b10001010;
   assign rom_data[1536]=8'b01000001;
   assign rom_data[1537]=8'b10001010;
   assign rom_data[1538]=8'b01000001;
   assign rom_data[1539]=8'b10001001;
   assign rom_data[1540]=8'b01000001;
   assign rom_data[1541]=8'b10001001;
   assign rom_data[1542]=8'b01000001;
   assign rom_data[1543]=8'b10001001;
   assign rom_data[1544]=8'b01000001;
   assign rom_data[1545]=8'b10001000;
   assign rom_data[1546]=8'b01000001;
   assign rom_data[1547]=8'b10001000;
   assign rom_data[1548]=8'b01000001;
   assign rom_data[1549]=8'b10000111;
   assign rom_data[1550]=8'b01000001;
   assign rom_data[1551]=8'b10000111;
   assign rom_data[1552]=8'b01000001;
   assign rom_data[1553]=8'b10000110;
   assign rom_data[1554]=8'b01000001;
   assign rom_data[1555]=8'b10000101;
   assign rom_data[1556]=8'b01000001;
   assign rom_data[1557]=8'b10000100;
   assign rom_data[1558]=8'b01000001;
   assign rom_data[1559]=8'b10000011;
   assign rom_data[1560]=8'b01000001;
   assign rom_data[1561]=8'b10000011;
   assign rom_data[1562]=8'b01000001;
   assign rom_data[1563]=8'b10000010;
   assign rom_data[1564]=8'b01000001;
   assign rom_data[1565]=8'b10000001;
   assign rom_data[1566]=8'b01000001;
   assign rom_data[1567]=8'b10000000;
   assign rom_data[1568]=8'b01000001;
   assign rom_data[1569]=8'b01111110;
   assign rom_data[1570]=8'b01000001;
   assign rom_data[1571]=8'b01111101;
   assign rom_data[1572]=8'b01000001;
   assign rom_data[1573]=8'b01111100;
   assign rom_data[1574]=8'b01000001;
   assign rom_data[1575]=8'b01111011;
   assign rom_data[1576]=8'b01000001;
   assign rom_data[1577]=8'b01111010;
   assign rom_data[1578]=8'b01000001;
   assign rom_data[1579]=8'b01111001;
   assign rom_data[1580]=8'b01000001;
   assign rom_data[1581]=8'b01110111;
   assign rom_data[1582]=8'b01000001;
   assign rom_data[1583]=8'b01110110;
   assign rom_data[1584]=8'b01000001;
   assign rom_data[1585]=8'b01110101;
   assign rom_data[1586]=8'b01000001;
   assign rom_data[1587]=8'b01110100;
   assign rom_data[1588]=8'b01000001;
   assign rom_data[1589]=8'b01110010;
   assign rom_data[1590]=8'b01000001;
   assign rom_data[1591]=8'b01110001;
   assign rom_data[1592]=8'b01000001;
   assign rom_data[1593]=8'b01110000;
   assign rom_data[1594]=8'b01000001;
   assign rom_data[1595]=8'b01101110;
   assign rom_data[1596]=8'b01000001;
   assign rom_data[1597]=8'b01101101;
   assign rom_data[1598]=8'b01000001;
   assign rom_data[1599]=8'b01101100;
   assign rom_data[1600]=8'b01000001;
   assign rom_data[1601]=8'b01101010;
   assign rom_data[1602]=8'b01000001;
   assign rom_data[1603]=8'b01101001;
   assign rom_data[1604]=8'b01000001;
   assign rom_data[1605]=8'b01100111;
   assign rom_data[1606]=8'b01000001;
   assign rom_data[1607]=8'b01100110;
   assign rom_data[1608]=8'b01000010;
   assign rom_data[1609]=8'b01100101;
   assign rom_data[1610]=8'b01000010;
   assign rom_data[1611]=8'b01100011;
   assign rom_data[1612]=8'b01000010;
   assign rom_data[1613]=8'b01100010;
   assign rom_data[1614]=8'b01000010;
   assign rom_data[1615]=8'b01100001;
   assign rom_data[1616]=8'b01000010;
   assign rom_data[1617]=8'b01011111;
   assign rom_data[1618]=8'b01000010;
   assign rom_data[1619]=8'b01011110;
   assign rom_data[1620]=8'b01000010;
   assign rom_data[1621]=8'b01011100;
   assign rom_data[1622]=8'b01000010;
   assign rom_data[1623]=8'b01011011;
   assign rom_data[1624]=8'b01000010;
   assign rom_data[1625]=8'b01011001;
   assign rom_data[1626]=8'b01000010;
   assign rom_data[1627]=8'b01011000;
   assign rom_data[1628]=8'b01000010;
   assign rom_data[1629]=8'b01010111;
   assign rom_data[1630]=8'b01000010;
   assign rom_data[1631]=8'b01010101;
   assign rom_data[1632]=8'b01000010;
   assign rom_data[1633]=8'b01010100;
   assign rom_data[1634]=8'b01000010;
   assign rom_data[1635]=8'b01010010;
   assign rom_data[1636]=8'b01000010;
   assign rom_data[1637]=8'b01010001;
   assign rom_data[1638]=8'b01000010;
   assign rom_data[1639]=8'b01010000;
   assign rom_data[1640]=8'b01000010;
   assign rom_data[1641]=8'b01001110;
   assign rom_data[1642]=8'b01000010;
   assign rom_data[1643]=8'b01001101;
   assign rom_data[1644]=8'b01000010;
   assign rom_data[1645]=8'b01001100;
   assign rom_data[1646]=8'b01000010;
   assign rom_data[1647]=8'b01001010;
   assign rom_data[1648]=8'b01000010;
   assign rom_data[1649]=8'b01001001;
   assign rom_data[1650]=8'b01000010;
   assign rom_data[1651]=8'b01001000;
   assign rom_data[1652]=8'b01000010;
   assign rom_data[1653]=8'b01000110;
   assign rom_data[1654]=8'b01000010;
   assign rom_data[1655]=8'b01000101;
   assign rom_data[1656]=8'b01000010;
   assign rom_data[1657]=8'b01000100;
   assign rom_data[1658]=8'b01000010;
   assign rom_data[1659]=8'b01000010;
   assign rom_data[1660]=8'b01000010;
   assign rom_data[1661]=8'b01000001;
   assign rom_data[1662]=8'b01000010;
   assign rom_data[1663]=8'b01000000;
   assign rom_data[1664]=8'b01000010;
   assign rom_data[1665]=8'b00111111;
   assign rom_data[1666]=8'b01000010;
   assign rom_data[1667]=8'b00111101;
   assign rom_data[1668]=8'b01000010;
   assign rom_data[1669]=8'b00111100;
   assign rom_data[1670]=8'b01000010;
   assign rom_data[1671]=8'b00111011;
   assign rom_data[1672]=8'b01000010;
   assign rom_data[1673]=8'b00111010;
   assign rom_data[1674]=8'b01000010;
   assign rom_data[1675]=8'b00111001;
   assign rom_data[1676]=8'b01000010;
   assign rom_data[1677]=8'b00111000;
   assign rom_data[1678]=8'b01000010;
   assign rom_data[1679]=8'b00110110;
   assign rom_data[1680]=8'b01000010;
   assign rom_data[1681]=8'b00110101;
   assign rom_data[1682]=8'b01000010;
   assign rom_data[1683]=8'b00110100;
   assign rom_data[1684]=8'b01000010;
   assign rom_data[1685]=8'b00110011;
   assign rom_data[1686]=8'b01000010;
   assign rom_data[1687]=8'b00110011;
   assign rom_data[1688]=8'b01000010;
   assign rom_data[1689]=8'b00110010;
   assign rom_data[1690]=8'b01000011;
   assign rom_data[1691]=8'b00110001;
   assign rom_data[1692]=8'b01000011;
   assign rom_data[1693]=8'b00110000;
   assign rom_data[1694]=8'b01000011;
   assign rom_data[1695]=8'b00101111;
   assign rom_data[1696]=8'b01000011;
   assign rom_data[1697]=8'b00101111;
   assign rom_data[1698]=8'b01000011;
   assign rom_data[1699]=8'b00101110;
   assign rom_data[1700]=8'b01000011;
   assign rom_data[1701]=8'b00101110;
   assign rom_data[1702]=8'b01000011;
   assign rom_data[1703]=8'b00101101;
   assign rom_data[1704]=8'b01000011;
   assign rom_data[1705]=8'b00101101;
   assign rom_data[1706]=8'b01000011;
   assign rom_data[1707]=8'b00101100;
   assign rom_data[1708]=8'b01000011;
   assign rom_data[1709]=8'b00101100;
   assign rom_data[1710]=8'b01000011;
   assign rom_data[1711]=8'b00101100;
   assign rom_data[1712]=8'b01000011;
   assign rom_data[1713]=8'b00101100;
   assign rom_data[1714]=8'b01000011;
   assign rom_data[1715]=8'b00101100;
   assign rom_data[1716]=8'b01000011;
   assign rom_data[1717]=8'b00101100;
   assign rom_data[1718]=8'b01000011;
   assign rom_data[1719]=8'b00101100;
   assign rom_data[1720]=8'b01000011;
   assign rom_data[1721]=8'b00101101;
   assign rom_data[1722]=8'b01000011;
   assign rom_data[1723]=8'b00101101;
   assign rom_data[1724]=8'b01000011;
   assign rom_data[1725]=8'b00101101;
   assign rom_data[1726]=8'b01000011;
   assign rom_data[1727]=8'b00101110;
   assign rom_data[1728]=8'b01000011;
   assign rom_data[1729]=8'b00101111;
   assign rom_data[1730]=8'b01000011;
   assign rom_data[1731]=8'b00101111;
   assign rom_data[1732]=8'b01000011;
   assign rom_data[1733]=8'b00110000;
   assign rom_data[1734]=8'b01000011;
   assign rom_data[1735]=8'b00110001;
   assign rom_data[1736]=8'b01000011;
   assign rom_data[1737]=8'b00110001;
   assign rom_data[1738]=8'b01000011;
   assign rom_data[1739]=8'b00110010;
   assign rom_data[1740]=8'b01000011;
   assign rom_data[1741]=8'b00110011;
   assign rom_data[1742]=8'b01000011;
   assign rom_data[1743]=8'b00110100;
   assign rom_data[1744]=8'b01000011;
   assign rom_data[1745]=8'b00110101;
   assign rom_data[1746]=8'b01000011;
   assign rom_data[1747]=8'b00110110;
   assign rom_data[1748]=8'b01000011;
   assign rom_data[1749]=8'b00110111;
   assign rom_data[1750]=8'b01000011;
   assign rom_data[1751]=8'b00111000;
   assign rom_data[1752]=8'b01000011;
   assign rom_data[1753]=8'b00111010;
   assign rom_data[1754]=8'b01000011;
   assign rom_data[1755]=8'b00111011;
   assign rom_data[1756]=8'b01000100;
   assign rom_data[1757]=8'b00111100;
   assign rom_data[1758]=8'b01000100;
   assign rom_data[1759]=8'b00111101;
   assign rom_data[1760]=8'b01000100;
   assign rom_data[1761]=8'b00111110;
   assign rom_data[1762]=8'b01000100;
   assign rom_data[1763]=8'b01000000;
   assign rom_data[1764]=8'b01000100;
   assign rom_data[1765]=8'b01000001;
   assign rom_data[1766]=8'b01000100;
   assign rom_data[1767]=8'b01000010;
   assign rom_data[1768]=8'b01000100;
   assign rom_data[1769]=8'b01000100;
   assign rom_data[1770]=8'b01000100;
   assign rom_data[1771]=8'b01000101;
   assign rom_data[1772]=8'b01000100;
   assign rom_data[1773]=8'b01000110;
   assign rom_data[1774]=8'b01000100;
   assign rom_data[1775]=8'b01000111;
   assign rom_data[1776]=8'b01000100;
   assign rom_data[1777]=8'b01001001;
   assign rom_data[1778]=8'b01000100;
   assign rom_data[1779]=8'b01001010;
   assign rom_data[1780]=8'b01000100;
   assign rom_data[1781]=8'b01001100;
   assign rom_data[1782]=8'b01000100;
   assign rom_data[1783]=8'b01001101;
   assign rom_data[1784]=8'b01000100;
   assign rom_data[1785]=8'b01001110;
   assign rom_data[1786]=8'b01000100;
   assign rom_data[1787]=8'b01010000;
   assign rom_data[1788]=8'b01000100;
   assign rom_data[1789]=8'b01010001;
   assign rom_data[1790]=8'b01000100;
   assign rom_data[1791]=8'b01010010;
   assign rom_data[1792]=8'b01000100;
   assign rom_data[1793]=8'b01010100;
   assign rom_data[1794]=8'b01000100;
   assign rom_data[1795]=8'b01010101;
   assign rom_data[1796]=8'b01000100;
   assign rom_data[1797]=8'b01010111;
   assign rom_data[1798]=8'b01000100;
   assign rom_data[1799]=8'b01011000;
   assign rom_data[1800]=8'b01000100;
   assign rom_data[1801]=8'b01011010;
   assign rom_data[1802]=8'b01000100;
   assign rom_data[1803]=8'b01011011;
   assign rom_data[1804]=8'b01000100;
   assign rom_data[1805]=8'b01011100;
   assign rom_data[1806]=8'b01000100;
   assign rom_data[1807]=8'b01011110;
   assign rom_data[1808]=8'b01000100;
   assign rom_data[1809]=8'b01011111;
   assign rom_data[1810]=8'b01000100;
   assign rom_data[1811]=8'b01100001;
   assign rom_data[1812]=8'b01000100;
   assign rom_data[1813]=8'b01100010;
   assign rom_data[1814]=8'b01000100;
   assign rom_data[1815]=8'b01100011;
   assign rom_data[1816]=8'b01000100;
   assign rom_data[1817]=8'b01100101;
   assign rom_data[1818]=8'b01000100;
   assign rom_data[1819]=8'b01100110;
   assign rom_data[1820]=8'b01000100;
   assign rom_data[1821]=8'b01100111;
   assign rom_data[1822]=8'b01000100;
   assign rom_data[1823]=8'b01101001;
   assign rom_data[1824]=8'b01000100;
   assign rom_data[1825]=8'b01101010;
   assign rom_data[1826]=8'b01000100;
   assign rom_data[1827]=8'b01101100;
   assign rom_data[1828]=8'b01000100;
   assign rom_data[1829]=8'b01101101;
   assign rom_data[1830]=8'b01000100;
   assign rom_data[1831]=8'b01101110;
   assign rom_data[1832]=8'b01000100;
   assign rom_data[1833]=8'b01110000;
   assign rom_data[1834]=8'b01000100;
   assign rom_data[1835]=8'b01110001;
   assign rom_data[1836]=8'b01000100;
   assign rom_data[1837]=8'b01110010;
   assign rom_data[1838]=8'b01000101;
   assign rom_data[1839]=8'b01110100;
   assign rom_data[1840]=8'b01000101;
   assign rom_data[1841]=8'b01110101;
   assign rom_data[1842]=8'b01000101;
   assign rom_data[1843]=8'b01110110;
   assign rom_data[1844]=8'b01000101;
   assign rom_data[1845]=8'b01110111;
   assign rom_data[1846]=8'b01000101;
   assign rom_data[1847]=8'b01111001;
   assign rom_data[1848]=8'b01000101;
   assign rom_data[1849]=8'b01111010;
   assign rom_data[1850]=8'b01000101;
   assign rom_data[1851]=8'b01111011;
   assign rom_data[1852]=8'b01000101;
   assign rom_data[1853]=8'b01111100;
   assign rom_data[1854]=8'b01000101;
   assign rom_data[1855]=8'b01111101;
   assign rom_data[1856]=8'b01000101;
   assign rom_data[1857]=8'b01111110;
   assign rom_data[1858]=8'b01000101;
   assign rom_data[1859]=8'b01111111;
   assign rom_data[1860]=8'b01000101;
   assign rom_data[1861]=8'b10000000;
   assign rom_data[1862]=8'b01000101;
   assign rom_data[1863]=8'b10000001;
   assign rom_data[1864]=8'b01000101;
   assign rom_data[1865]=8'b10000010;
   assign rom_data[1866]=8'b01000101;
   assign rom_data[1867]=8'b10000011;
   assign rom_data[1868]=8'b01000101;
   assign rom_data[1869]=8'b10000100;
   assign rom_data[1870]=8'b01000101;
   assign rom_data[1871]=8'b10000101;
   assign rom_data[1872]=8'b01000101;
   assign rom_data[1873]=8'b10000110;
   assign rom_data[1874]=8'b01000101;
   assign rom_data[1875]=8'b10000110;
   assign rom_data[1876]=8'b01000101;
   assign rom_data[1877]=8'b10000111;
   assign rom_data[1878]=8'b01000101;
   assign rom_data[1879]=8'b10001000;
   assign rom_data[1880]=8'b01000101;
   assign rom_data[1881]=8'b10001000;
   assign rom_data[1882]=8'b01000101;
   assign rom_data[1883]=8'b10001001;
   assign rom_data[1884]=8'b01000101;
   assign rom_data[1885]=8'b10001001;
   assign rom_data[1886]=8'b01000101;
   assign rom_data[1887]=8'b10001001;
   assign rom_data[1888]=8'b01000101;
   assign rom_data[1889]=8'b10001010;
   assign rom_data[1890]=8'b01000101;
   assign rom_data[1891]=8'b10001010;
   assign rom_data[1892]=8'b01000101;
   assign rom_data[1893]=8'b10001010;
   assign rom_data[1894]=8'b01000101;
   assign rom_data[1895]=8'b10001010;
   assign rom_data[1896]=8'b01000101;
   assign rom_data[1897]=8'b10001010;
   assign rom_data[1898]=8'b01000101;
   assign rom_data[1899]=8'b10001001;
   assign rom_data[1900]=8'b01000101;
   assign rom_data[1901]=8'b10001001;
   assign rom_data[1902]=8'b01000101;
   assign rom_data[1903]=8'b10001001;
   assign rom_data[1904]=8'b01000101;
   assign rom_data[1905]=8'b10001000;
   assign rom_data[1906]=8'b01000101;
   assign rom_data[1907]=8'b10001000;
   assign rom_data[1908]=8'b01000110;
   assign rom_data[1909]=8'b10000111;
   assign rom_data[1910]=8'b01000110;
   assign rom_data[1911]=8'b10000111;
   assign rom_data[1912]=8'b01000110;
   assign rom_data[1913]=8'b10000110;
   assign rom_data[1914]=8'b01000110;
   assign rom_data[1915]=8'b10000101;
   assign rom_data[1916]=8'b01000110;
   assign rom_data[1917]=8'b10000100;
   assign rom_data[1918]=8'b01000110;
   assign rom_data[1919]=8'b10000011;
   assign rom_data[1920]=8'b01000110;
   assign rom_data[1921]=8'b10000011;
   assign rom_data[1922]=8'b01000110;
   assign rom_data[1923]=8'b10000010;
   assign rom_data[1924]=8'b01000110;
   assign rom_data[1925]=8'b10000001;
   assign rom_data[1926]=8'b01000110;
   assign rom_data[1927]=8'b10000000;
   assign rom_data[1928]=8'b01000110;
   assign rom_data[1929]=8'b01111110;
   assign rom_data[1930]=8'b01000110;
   assign rom_data[1931]=8'b01111101;
   assign rom_data[1932]=8'b01000110;
   assign rom_data[1933]=8'b01111100;
   assign rom_data[1934]=8'b01000110;
   assign rom_data[1935]=8'b01111011;
   assign rom_data[1936]=8'b01000110;
   assign rom_data[1937]=8'b01111010;
   assign rom_data[1938]=8'b01000110;
   assign rom_data[1939]=8'b01111001;
   assign rom_data[1940]=8'b01000110;
   assign rom_data[1941]=8'b01110111;
   assign rom_data[1942]=8'b01000110;
   assign rom_data[1943]=8'b01110110;
   assign rom_data[1944]=8'b01000110;
   assign rom_data[1945]=8'b01110101;
   assign rom_data[1946]=8'b01000110;
   assign rom_data[1947]=8'b01110100;
   assign rom_data[1948]=8'b01000110;
   assign rom_data[1949]=8'b01110010;
   assign rom_data[1950]=8'b01000110;
   assign rom_data[1951]=8'b01110001;
   assign rom_data[1952]=8'b01000110;
   assign rom_data[1953]=8'b01110000;
   assign rom_data[1954]=8'b01000110;
   assign rom_data[1955]=8'b01101110;
   assign rom_data[1956]=8'b01000110;
   assign rom_data[1957]=8'b01101101;
   assign rom_data[1958]=8'b01000110;
   assign rom_data[1959]=8'b01101100;
   assign rom_data[1960]=8'b01000110;
   assign rom_data[1961]=8'b01101010;
   assign rom_data[1962]=8'b01000110;
   assign rom_data[1963]=8'b01101001;
   assign rom_data[1964]=8'b01000110;
   assign rom_data[1965]=8'b01100111;
   assign rom_data[1966]=8'b01000110;
   assign rom_data[1967]=8'b01100110;
   assign rom_data[1968]=8'b01000110;
   assign rom_data[1969]=8'b01100101;
   assign rom_data[1970]=8'b01000110;
   assign rom_data[1971]=8'b01100011;
   assign rom_data[1972]=8'b01000110;
   assign rom_data[1973]=8'b01100010;
   assign rom_data[1974]=8'b01000110;
   assign rom_data[1975]=8'b01100001;
   assign rom_data[1976]=8'b01000110;
   assign rom_data[1977]=8'b01011111;
   assign rom_data[1978]=8'b01000110;
   assign rom_data[1979]=8'b01011110;
   assign rom_data[1980]=8'b01000110;
   assign rom_data[1981]=8'b01011100;
   assign rom_data[1982]=8'b01000110;
   assign rom_data[1983]=8'b01011011;
   assign rom_data[1984]=8'b01000111;
   assign rom_data[1985]=8'b01011001;
   assign rom_data[1986]=8'b01000111;
   assign rom_data[1987]=8'b01011000;
   assign rom_data[1988]=8'b01000111;
   assign rom_data[1989]=8'b01010111;
   assign rom_data[1990]=8'b01000111;
   assign rom_data[1991]=8'b01010101;
   assign rom_data[1992]=8'b01000111;
   assign rom_data[1993]=8'b01010100;
   assign rom_data[1994]=8'b01000111;
   assign rom_data[1995]=8'b01010010;
   assign rom_data[1996]=8'b01000111;
   assign rom_data[1997]=8'b01010001;
   assign rom_data[1998]=8'b01000111;
   assign rom_data[1999]=8'b01010000;
   assign rom_data[2000]=8'b01000111;
   assign rom_data[2001]=8'b01001110;
   assign rom_data[2002]=8'b01000111;
   assign rom_data[2003]=8'b01001101;
   assign rom_data[2004]=8'b01000111;
   assign rom_data[2005]=8'b01001100;
   assign rom_data[2006]=8'b01000111;
   assign rom_data[2007]=8'b01001010;
   assign rom_data[2008]=8'b01000111;
   assign rom_data[2009]=8'b01001001;
   assign rom_data[2010]=8'b01000111;
   assign rom_data[2011]=8'b01001000;
   assign rom_data[2012]=8'b01000111;
   assign rom_data[2013]=8'b01000110;
   assign rom_data[2014]=8'b01000111;
   assign rom_data[2015]=8'b01000101;
   assign rom_data[2016]=8'b01000111;
   assign rom_data[2017]=8'b01000100;
   assign rom_data[2018]=8'b01000111;
   assign rom_data[2019]=8'b01000010;
   assign rom_data[2020]=8'b01000111;
   assign rom_data[2021]=8'b01000001;
   assign rom_data[2022]=8'b01000111;
   assign rom_data[2023]=8'b01000000;
   assign rom_data[2024]=8'b01000111;
   assign rom_data[2025]=8'b00111111;
   assign rom_data[2026]=8'b01000111;
   assign rom_data[2027]=8'b00111101;
   assign rom_data[2028]=8'b01000111;
   assign rom_data[2029]=8'b00111100;
   assign rom_data[2030]=8'b01000111;
   assign rom_data[2031]=8'b00111011;
   assign rom_data[2032]=8'b01000111;
   assign rom_data[2033]=8'b00111010;
   assign rom_data[2034]=8'b01000111;
   assign rom_data[2035]=8'b00111001;
   assign rom_data[2036]=8'b01000111;
   assign rom_data[2037]=8'b00111000;
   assign rom_data[2038]=8'b01000111;
   assign rom_data[2039]=8'b00110110;
   assign rom_data[2040]=8'b01000111;
   assign rom_data[2041]=8'b00110101;
   assign rom_data[2042]=8'b01000111;
   assign rom_data[2043]=8'b00110100;
   assign rom_data[2044]=8'b01000111;
   assign rom_data[2045]=8'b00110011;
   assign rom_data[2046]=8'b01000111;
   assign rom_data[2047]=8'b00110011;
   assign rom_data[2048]=8'b01000111;
   assign rom_data[2049]=8'b00110010;
   assign rom_data[2050]=8'b01000111;
   assign rom_data[2051]=8'b00110001;
   assign rom_data[2052]=8'b01000111;
   assign rom_data[2053]=8'b00110000;
   assign rom_data[2054]=8'b01000111;
   assign rom_data[2055]=8'b00101111;
   assign rom_data[2056]=8'b01000111;
   assign rom_data[2057]=8'b00101111;
   assign rom_data[2058]=8'b01000111;
   assign rom_data[2059]=8'b00101110;
   assign rom_data[2060]=8'b01000111;
   assign rom_data[2061]=8'b00101110;
   assign rom_data[2062]=8'b01001000;
   assign rom_data[2063]=8'b00101101;
   assign rom_data[2064]=8'b01001000;
   assign rom_data[2065]=8'b00101101;
   assign rom_data[2066]=8'b01001000;
   assign rom_data[2067]=8'b00101100;
   assign rom_data[2068]=8'b01001000;
   assign rom_data[2069]=8'b00101100;
   assign rom_data[2070]=8'b01001000;
   assign rom_data[2071]=8'b00101100;
   assign rom_data[2072]=8'b01001000;
   assign rom_data[2073]=8'b00101100;
   assign rom_data[2074]=8'b01001000;
   assign rom_data[2075]=8'b00101100;
   assign rom_data[2076]=8'b01001000;
   assign rom_data[2077]=8'b00101100;
   assign rom_data[2078]=8'b01001000;
   assign rom_data[2079]=8'b00101100;
   assign rom_data[2080]=8'b01001000;
   assign rom_data[2081]=8'b00101101;
   assign rom_data[2082]=8'b01001000;
   assign rom_data[2083]=8'b00101101;
   assign rom_data[2084]=8'b01001000;
   assign rom_data[2085]=8'b00101101;
   assign rom_data[2086]=8'b01001000;
   assign rom_data[2087]=8'b00101110;
   assign rom_data[2088]=8'b01001000;
   assign rom_data[2089]=8'b00101111;
   assign rom_data[2090]=8'b01001000;
   assign rom_data[2091]=8'b00101111;
   assign rom_data[2092]=8'b01001000;
   assign rom_data[2093]=8'b00110000;
   assign rom_data[2094]=8'b01001000;
   assign rom_data[2095]=8'b00110001;
   assign rom_data[2096]=8'b01001000;
   assign rom_data[2097]=8'b00110001;
   assign rom_data[2098]=8'b01001000;
   assign rom_data[2099]=8'b00110010;
   assign rom_data[2100]=8'b01001000;
   assign rom_data[2101]=8'b00110011;
   assign rom_data[2102]=8'b01001000;
   assign rom_data[2103]=8'b00110100;
   assign rom_data[2104]=8'b01001000;
   assign rom_data[2105]=8'b00110101;
   assign rom_data[2106]=8'b01001000;
   assign rom_data[2107]=8'b00110110;
   assign rom_data[2108]=8'b01001000;
   assign rom_data[2109]=8'b00110111;
   assign rom_data[2110]=8'b01001000;
   assign rom_data[2111]=8'b00111000;
   assign rom_data[2112]=8'b01001000;
   assign rom_data[2113]=8'b00111010;
   assign rom_data[2114]=8'b01001000;
   assign rom_data[2115]=8'b00111011;
   assign rom_data[2116]=8'b01001000;
   assign rom_data[2117]=8'b00111100;
   assign rom_data[2118]=8'b01001000;
   assign rom_data[2119]=8'b00111101;
   assign rom_data[2120]=8'b01001000;
   assign rom_data[2121]=8'b00111110;
   assign rom_data[2122]=8'b01001000;
   assign rom_data[2123]=8'b01000000;
   assign rom_data[2124]=8'b01001000;
   assign rom_data[2125]=8'b01000001;
   assign rom_data[2126]=8'b01001000;
   assign rom_data[2127]=8'b01000010;
   assign rom_data[2128]=8'b01001000;
   assign rom_data[2129]=8'b01000100;
   assign rom_data[2130]=8'b01001001;
   assign rom_data[2131]=8'b01000101;
   assign rom_data[2132]=8'b01001001;
   assign rom_data[2133]=8'b01000110;
   assign rom_data[2134]=8'b01001001;
   assign rom_data[2135]=8'b01000111;
   assign rom_data[2136]=8'b01001001;
   assign rom_data[2137]=8'b01001001;
   assign rom_data[2138]=8'b01001001;
   assign rom_data[2139]=8'b01001010;
   assign rom_data[2140]=8'b01001001;
   assign rom_data[2141]=8'b01001100;
   assign rom_data[2142]=8'b01001001;
   assign rom_data[2143]=8'b01001101;
   assign rom_data[2144]=8'b01001001;
   assign rom_data[2145]=8'b01001110;
   assign rom_data[2146]=8'b01001001;
   assign rom_data[2147]=8'b01010000;
   assign rom_data[2148]=8'b01001001;
   assign rom_data[2149]=8'b01010001;
   assign rom_data[2150]=8'b01001001;
   assign rom_data[2151]=8'b01010010;
   assign rom_data[2152]=8'b01001001;
   assign rom_data[2153]=8'b01010100;
   assign rom_data[2154]=8'b01001001;
   assign rom_data[2155]=8'b01010101;
   assign rom_data[2156]=8'b01001001;
   assign rom_data[2157]=8'b01010111;
   assign rom_data[2158]=8'b01001001;
   assign rom_data[2159]=8'b01011000;
   assign rom_data[2160]=8'b01001001;
   assign rom_data[2161]=8'b01011010;
   assign rom_data[2162]=8'b01001001;
   assign rom_data[2163]=8'b01011011;
   assign rom_data[2164]=8'b01001001;
   assign rom_data[2165]=8'b01011100;
   assign rom_data[2166]=8'b01001001;
   assign rom_data[2167]=8'b01011110;
   assign rom_data[2168]=8'b01001001;
   assign rom_data[2169]=8'b01011111;
   assign rom_data[2170]=8'b01001001;
   assign rom_data[2171]=8'b01100001;
   assign rom_data[2172]=8'b01001001;
   assign rom_data[2173]=8'b01100010;
   assign rom_data[2174]=8'b01001001;
   assign rom_data[2175]=8'b01100011;
   assign rom_data[2176]=8'b01001001;
   assign rom_data[2177]=8'b01100101;
   assign rom_data[2178]=8'b01001001;
   assign rom_data[2179]=8'b01100110;
   assign rom_data[2180]=8'b01001001;
   assign rom_data[2181]=8'b01100111;
   assign rom_data[2182]=8'b01001001;
   assign rom_data[2183]=8'b01101001;
   assign rom_data[2184]=8'b01001001;
   assign rom_data[2185]=8'b01101010;
   assign rom_data[2186]=8'b01001001;
   assign rom_data[2187]=8'b01101100;
   assign rom_data[2188]=8'b01001001;
   assign rom_data[2189]=8'b01101101;
   assign rom_data[2190]=8'b01001001;
   assign rom_data[2191]=8'b01101110;
   assign rom_data[2192]=8'b01001001;
   assign rom_data[2193]=8'b01110000;
   assign rom_data[2194]=8'b01001001;
   assign rom_data[2195]=8'b01110001;
   assign rom_data[2196]=8'b01001001;
   assign rom_data[2197]=8'b01110010;
   assign rom_data[2198]=8'b01001001;
   assign rom_data[2199]=8'b01110100;
   assign rom_data[2200]=8'b01001001;
   assign rom_data[2201]=8'b01110101;
   assign rom_data[2202]=8'b01001001;
   assign rom_data[2203]=8'b01110110;
   assign rom_data[2204]=8'b01001001;
   assign rom_data[2205]=8'b01110111;
   assign rom_data[2206]=8'b01001001;
   assign rom_data[2207]=8'b01111001;
   assign rom_data[2208]=8'b01001001;
   assign rom_data[2209]=8'b01111010;
   assign rom_data[2210]=8'b01001001;
   assign rom_data[2211]=8'b01111011;
   assign rom_data[2212]=8'b01001001;
   assign rom_data[2213]=8'b01111100;
   assign rom_data[2214]=8'b01001010;
   assign rom_data[2215]=8'b01111101;
   assign rom_data[2216]=8'b01001010;
   assign rom_data[2217]=8'b01111110;
   assign rom_data[2218]=8'b01001010;
   assign rom_data[2219]=8'b01111111;
   assign rom_data[2220]=8'b01001010;
   assign rom_data[2221]=8'b10000000;
   assign rom_data[2222]=8'b01001010;
   assign rom_data[2223]=8'b10000001;
   assign rom_data[2224]=8'b01001010;
   assign rom_data[2225]=8'b10000010;
   assign rom_data[2226]=8'b01001010;
   assign rom_data[2227]=8'b10000011;
   assign rom_data[2228]=8'b01001010;
   assign rom_data[2229]=8'b10000100;
   assign rom_data[2230]=8'b01001010;
   assign rom_data[2231]=8'b10000101;
   assign rom_data[2232]=8'b01001010;
   assign rom_data[2233]=8'b10000110;
   assign rom_data[2234]=8'b01001010;
   assign rom_data[2235]=8'b10000110;
   assign rom_data[2236]=8'b01001010;
   assign rom_data[2237]=8'b10000111;
   assign rom_data[2238]=8'b01001010;
   assign rom_data[2239]=8'b10001000;
   assign rom_data[2240]=8'b01001010;
   assign rom_data[2241]=8'b10001000;
   assign rom_data[2242]=8'b01001010;
   assign rom_data[2243]=8'b10001001;
   assign rom_data[2244]=8'b01001010;
   assign rom_data[2245]=8'b10001001;
   assign rom_data[2246]=8'b01001010;
   assign rom_data[2247]=8'b10001001;
   assign rom_data[2248]=8'b01001010;
   assign rom_data[2249]=8'b10001010;
   assign rom_data[2250]=8'b01001010;
   assign rom_data[2251]=8'b10001010;
   assign rom_data[2252]=8'b01001010;
   assign rom_data[2253]=8'b10001010;
   assign rom_data[2254]=8'b01001010;
   assign rom_data[2255]=8'b10001010;
   assign rom_data[2256]=8'b01001010;
   assign rom_data[2257]=8'b10001010;
   assign rom_data[2258]=8'b01001010;
   assign rom_data[2259]=8'b10001001;
   assign rom_data[2260]=8'b01001010;
   assign rom_data[2261]=8'b10001001;
   assign rom_data[2262]=8'b01001010;
   assign rom_data[2263]=8'b10001001;
   assign rom_data[2264]=8'b01001010;
   assign rom_data[2265]=8'b10001000;
   assign rom_data[2266]=8'b01001010;
   assign rom_data[2267]=8'b10001000;
   assign rom_data[2268]=8'b01001010;
   assign rom_data[2269]=8'b10000111;
   assign rom_data[2270]=8'b01001010;
   assign rom_data[2271]=8'b10000111;
   assign rom_data[2272]=8'b01001010;
   assign rom_data[2273]=8'b10000110;
   assign rom_data[2274]=8'b01001010;
   assign rom_data[2275]=8'b10000101;
   assign rom_data[2276]=8'b01001010;
   assign rom_data[2277]=8'b10000100;
   assign rom_data[2278]=8'b01001010;
   assign rom_data[2279]=8'b10000011;
   assign rom_data[2280]=8'b01001011;
   assign rom_data[2281]=8'b10000011;
   assign rom_data[2282]=8'b01001011;
   assign rom_data[2283]=8'b10000010;
   assign rom_data[2284]=8'b01001011;
   assign rom_data[2285]=8'b10000001;
   assign rom_data[2286]=8'b01001011;
   assign rom_data[2287]=8'b10000000;
   assign rom_data[2288]=8'b01001011;
   assign rom_data[2289]=8'b01111110;
   assign rom_data[2290]=8'b01001011;
   assign rom_data[2291]=8'b01111101;
   assign rom_data[2292]=8'b01001011;
   assign rom_data[2293]=8'b01111100;
   assign rom_data[2294]=8'b01001011;
   assign rom_data[2295]=8'b01111011;
   assign rom_data[2296]=8'b01001011;
   assign rom_data[2297]=8'b01111010;
   assign rom_data[2298]=8'b01001011;
   assign rom_data[2299]=8'b01111001;
   assign rom_data[2300]=8'b01001011;
   assign rom_data[2301]=8'b01110111;
   assign rom_data[2302]=8'b01001011;
   assign rom_data[2303]=8'b01110110;
   assign rom_data[2304]=8'b01001011;
   assign rom_data[2305]=8'b01110101;
   assign rom_data[2306]=8'b01001011;
   assign rom_data[2307]=8'b01110100;
   assign rom_data[2308]=8'b01001011;
   assign rom_data[2309]=8'b01110010;
   assign rom_data[2310]=8'b01001011;
   assign rom_data[2311]=8'b01110001;
   assign rom_data[2312]=8'b01001011;
   assign rom_data[2313]=8'b01110000;
   assign rom_data[2314]=8'b01001011;
   assign rom_data[2315]=8'b01101110;
   assign rom_data[2316]=8'b01001011;
   assign rom_data[2317]=8'b01101101;
   assign rom_data[2318]=8'b01001011;
   assign rom_data[2319]=8'b01101100;
   assign rom_data[2320]=8'b01001011;
   assign rom_data[2321]=8'b01101010;
   assign rom_data[2322]=8'b01001011;
   assign rom_data[2323]=8'b01101001;
   assign rom_data[2324]=8'b01001011;
   assign rom_data[2325]=8'b01100111;
   assign rom_data[2326]=8'b01001011;
   assign rom_data[2327]=8'b01100110;
   assign rom_data[2328]=8'b01001011;
   assign rom_data[2329]=8'b01100101;
   assign rom_data[2330]=8'b01001011;
   assign rom_data[2331]=8'b01100011;
   assign rom_data[2332]=8'b01001011;
   assign rom_data[2333]=8'b01100010;
   assign rom_data[2334]=8'b01001011;
   assign rom_data[2335]=8'b01100001;
   assign rom_data[2336]=8'b01001011;
   assign rom_data[2337]=8'b01011111;
   assign rom_data[2338]=8'b01001011;
   assign rom_data[2339]=8'b01011110;
   assign rom_data[2340]=8'b01001011;
   assign rom_data[2341]=8'b01011100;
   assign rom_data[2342]=8'b01001011;
   assign rom_data[2343]=8'b01011011;
   assign rom_data[2344]=8'b01001011;
   assign rom_data[2345]=8'b01011001;
   assign rom_data[2346]=8'b01001011;
   assign rom_data[2347]=8'b01011000;
   assign rom_data[2348]=8'b01001011;
   assign rom_data[2349]=8'b01010111;
   assign rom_data[2350]=8'b01001011;
   assign rom_data[2351]=8'b01010101;
   assign rom_data[2352]=8'b01001011;
   assign rom_data[2353]=8'b01010100;
   assign rom_data[2354]=8'b01001011;
   assign rom_data[2355]=8'b01010010;
   assign rom_data[2356]=8'b01001011;
   assign rom_data[2357]=8'b01010001;
   assign rom_data[2358]=8'b01001011;
   assign rom_data[2359]=8'b01010000;
   assign rom_data[2360]=8'b01001011;
   assign rom_data[2361]=8'b01001110;
   assign rom_data[2362]=8'b01001100;
   assign rom_data[2363]=8'b01001101;
   assign rom_data[2364]=8'b01001100;
   assign rom_data[2365]=8'b01001100;
   assign rom_data[2366]=8'b01001100;
   assign rom_data[2367]=8'b01001010;
   assign rom_data[2368]=8'b01001100;
   assign rom_data[2369]=8'b01001001;
   assign rom_data[2370]=8'b01001100;
   assign rom_data[2371]=8'b01001000;
   assign rom_data[2372]=8'b01001100;
   assign rom_data[2373]=8'b01000110;
   assign rom_data[2374]=8'b01001100;
   assign rom_data[2375]=8'b01000101;
   assign rom_data[2376]=8'b01001100;
   assign rom_data[2377]=8'b01000100;
   assign rom_data[2378]=8'b01001100;
   assign rom_data[2379]=8'b01000010;
   assign rom_data[2380]=8'b01001100;
   assign rom_data[2381]=8'b01000001;
   assign rom_data[2382]=8'b01001100;
   assign rom_data[2383]=8'b01000000;
   assign rom_data[2384]=8'b01001100;
   assign rom_data[2385]=8'b00111111;
   assign rom_data[2386]=8'b01001100;
   assign rom_data[2387]=8'b00111101;
   assign rom_data[2388]=8'b01001100;
   assign rom_data[2389]=8'b00111100;
   assign rom_data[2390]=8'b01001100;
   assign rom_data[2391]=8'b00111011;
   assign rom_data[2392]=8'b01001100;
   assign rom_data[2393]=8'b00111010;
   assign rom_data[2394]=8'b01001100;
   assign rom_data[2395]=8'b00111001;
   assign rom_data[2396]=8'b01001100;
   assign rom_data[2397]=8'b00111000;
   assign rom_data[2398]=8'b01001100;
   assign rom_data[2399]=8'b00110110;
   assign rom_data[2400]=8'b01001100;
   assign rom_data[2401]=8'b00110101;
   assign rom_data[2402]=8'b01001100;
   assign rom_data[2403]=8'b00110100;
   assign rom_data[2404]=8'b01001100;
   assign rom_data[2405]=8'b00110011;
   assign rom_data[2406]=8'b01001100;
   assign rom_data[2407]=8'b00110011;
   assign rom_data[2408]=8'b01001100;
   assign rom_data[2409]=8'b00110010;
   assign rom_data[2410]=8'b01001100;
   assign rom_data[2411]=8'b00110001;
   assign rom_data[2412]=8'b01001100;
   assign rom_data[2413]=8'b00110000;
   assign rom_data[2414]=8'b01001100;
   assign rom_data[2415]=8'b00101111;
   assign rom_data[2416]=8'b01001100;
   assign rom_data[2417]=8'b00101111;
   assign rom_data[2418]=8'b01001100;
   assign rom_data[2419]=8'b00101110;
   assign rom_data[2420]=8'b01001100;
   assign rom_data[2421]=8'b00101110;
   assign rom_data[2422]=8'b01001100;
   assign rom_data[2423]=8'b00101101;
   assign rom_data[2424]=8'b01001100;
   assign rom_data[2425]=8'b00101101;
   assign rom_data[2426]=8'b01001100;
   assign rom_data[2427]=8'b00101100;
   assign rom_data[2428]=8'b01001100;
   assign rom_data[2429]=8'b00101100;
   assign rom_data[2430]=8'b01001100;
   assign rom_data[2431]=8'b00101100;
   assign rom_data[2432]=8'b01001100;
   assign rom_data[2433]=8'b00101100;
   assign rom_data[2434]=8'b01001101;
   assign rom_data[2435]=8'b00101100;
   assign rom_data[2436]=8'b01001101;
   assign rom_data[2437]=8'b00101100;
   assign rom_data[2438]=8'b01001101;
   assign rom_data[2439]=8'b00101100;
   assign rom_data[2440]=8'b01001101;
   assign rom_data[2441]=8'b00101101;
   assign rom_data[2442]=8'b01001101;
   assign rom_data[2443]=8'b00101101;
   assign rom_data[2444]=8'b01001101;
   assign rom_data[2445]=8'b00101101;
   assign rom_data[2446]=8'b01001101;
   assign rom_data[2447]=8'b00101110;
   assign rom_data[2448]=8'b01001101;
   assign rom_data[2449]=8'b00101111;
   assign rom_data[2450]=8'b01001101;
   assign rom_data[2451]=8'b00101111;
   assign rom_data[2452]=8'b01001101;
   assign rom_data[2453]=8'b00110000;
   assign rom_data[2454]=8'b01001101;
   assign rom_data[2455]=8'b00110001;
   assign rom_data[2456]=8'b01001101;
   assign rom_data[2457]=8'b00110001;
   assign rom_data[2458]=8'b01001101;
   assign rom_data[2459]=8'b00110010;
   assign rom_data[2460]=8'b01001101;
   assign rom_data[2461]=8'b00110011;
   assign rom_data[2462]=8'b01001101;
   assign rom_data[2463]=8'b00110100;
   assign rom_data[2464]=8'b01001101;
   assign rom_data[2465]=8'b00110101;
   assign rom_data[2466]=8'b01001101;
   assign rom_data[2467]=8'b00110110;
   assign rom_data[2468]=8'b01001101;
   assign rom_data[2469]=8'b00110111;
   assign rom_data[2470]=8'b01001101;
   assign rom_data[2471]=8'b00111000;
   assign rom_data[2472]=8'b01001101;
   assign rom_data[2473]=8'b00111010;
   assign rom_data[2474]=8'b01001101;
   assign rom_data[2475]=8'b00111011;
   assign rom_data[2476]=8'b01001101;
   assign rom_data[2477]=8'b00111100;
   assign rom_data[2478]=8'b01001101;
   assign rom_data[2479]=8'b00111101;
   assign rom_data[2480]=8'b01001101;
   assign rom_data[2481]=8'b00111110;
   assign rom_data[2482]=8'b01001101;
   assign rom_data[2483]=8'b01000000;
   assign rom_data[2484]=8'b01001101;
   assign rom_data[2485]=8'b01000001;
   assign rom_data[2486]=8'b01001101;
   assign rom_data[2487]=8'b01000010;
   assign rom_data[2488]=8'b01001101;
   assign rom_data[2489]=8'b01000100;
   assign rom_data[2490]=8'b01001101;
   assign rom_data[2491]=8'b01000101;
   assign rom_data[2492]=8'b01001101;
   assign rom_data[2493]=8'b01000110;
   assign rom_data[2494]=8'b01001101;
   assign rom_data[2495]=8'b01000111;
   assign rom_data[2496]=8'b01001101;
   assign rom_data[2497]=8'b01001001;
   assign rom_data[2498]=8'b01001101;
   assign rom_data[2499]=8'b01001010;
   assign rom_data[2500]=8'b01001101;
   assign rom_data[2501]=8'b01001100;
   assign rom_data[2502]=8'b01001101;
   assign rom_data[2503]=8'b01001101;
   assign rom_data[2504]=8'b01001101;
   assign rom_data[2505]=8'b01001110;
   assign rom_data[2506]=8'b01001110;
   assign rom_data[2507]=8'b01010000;
   assign rom_data[2508]=8'b01001110;
   assign rom_data[2509]=8'b01010001;
   assign rom_data[2510]=8'b01001110;
   assign rom_data[2511]=8'b01010010;
   assign rom_data[2512]=8'b01001110;
   assign rom_data[2513]=8'b01010100;
   assign rom_data[2514]=8'b01001110;
   assign rom_data[2515]=8'b01010101;
   assign rom_data[2516]=8'b01001110;
   assign rom_data[2517]=8'b01010111;
   assign rom_data[2518]=8'b01001110;
   assign rom_data[2519]=8'b01011000;
   assign rom_data[2520]=8'b01001110;
   assign rom_data[2521]=8'b01011010;
   assign rom_data[2522]=8'b01001110;
   assign rom_data[2523]=8'b01011011;
   assign rom_data[2524]=8'b01001110;
   assign rom_data[2525]=8'b01011100;
   assign rom_data[2526]=8'b01001110;
   assign rom_data[2527]=8'b01011110;
   assign rom_data[2528]=8'b01001110;
   assign rom_data[2529]=8'b01011111;
   assign rom_data[2530]=8'b01001110;
   assign rom_data[2531]=8'b01100001;
   assign rom_data[2532]=8'b01001110;
   assign rom_data[2533]=8'b01100010;
   assign rom_data[2534]=8'b01001110;
   assign rom_data[2535]=8'b01100011;
   assign rom_data[2536]=8'b01001110;
   assign rom_data[2537]=8'b01100101;
   assign rom_data[2538]=8'b01001110;
   assign rom_data[2539]=8'b01100110;
   assign rom_data[2540]=8'b01001110;
   assign rom_data[2541]=8'b01100111;
   assign rom_data[2542]=8'b01001110;
   assign rom_data[2543]=8'b01101001;
   assign rom_data[2544]=8'b01001110;
   assign rom_data[2545]=8'b01101010;
   assign rom_data[2546]=8'b01001110;
   assign rom_data[2547]=8'b01101100;
   assign rom_data[2548]=8'b01001110;
   assign rom_data[2549]=8'b01101101;
   assign rom_data[2550]=8'b01001110;
   assign rom_data[2551]=8'b01101110;
   assign rom_data[2552]=8'b01001110;
   assign rom_data[2553]=8'b01110000;
   assign rom_data[2554]=8'b01001110;
   assign rom_data[2555]=8'b01110001;
   assign rom_data[2556]=8'b01001110;
   assign rom_data[2557]=8'b01110010;
   assign rom_data[2558]=8'b01001110;
   assign rom_data[2559]=8'b01110100;
   assign rom_data[2560]=8'b01001110;
   assign rom_data[2561]=8'b01110101;
   assign rom_data[2562]=8'b01001110;
   assign rom_data[2563]=8'b01110110;
   assign rom_data[2564]=8'b01001110;
   assign rom_data[2565]=8'b01110111;
   assign rom_data[2566]=8'b01001110;
   assign rom_data[2567]=8'b01111001;
   assign rom_data[2568]=8'b01001110;
   assign rom_data[2569]=8'b01111010;
   assign rom_data[2570]=8'b01001110;
   assign rom_data[2571]=8'b01111011;
   assign rom_data[2572]=8'b01001110;
   assign rom_data[2573]=8'b01111100;
   assign rom_data[2574]=8'b01001110;
   assign rom_data[2575]=8'b01111101;
   assign rom_data[2576]=8'b01001110;
   assign rom_data[2577]=8'b01111110;
   assign rom_data[2578]=8'b01001110;
   assign rom_data[2579]=8'b01111111;
   assign rom_data[2580]=8'b01001110;
   assign rom_data[2581]=8'b10000000;
   assign rom_data[2582]=8'b01001110;
   assign rom_data[2583]=8'b10000001;
   assign rom_data[2584]=8'b01001110;
   assign rom_data[2585]=8'b10000010;
   assign rom_data[2586]=8'b01001110;
   assign rom_data[2587]=8'b10000011;
   assign rom_data[2588]=8'b01001111;
   assign rom_data[2589]=8'b10000100;
   assign rom_data[2590]=8'b01001111;
   assign rom_data[2591]=8'b10000101;
   assign rom_data[2592]=8'b01001111;
   assign rom_data[2593]=8'b10000110;
   assign rom_data[2594]=8'b01001111;
   assign rom_data[2595]=8'b10000110;
   assign rom_data[2596]=8'b01001111;
   assign rom_data[2597]=8'b10000111;
   assign rom_data[2598]=8'b01001111;
   assign rom_data[2599]=8'b10001000;
   assign rom_data[2600]=8'b01001111;
   assign rom_data[2601]=8'b10001000;
   assign rom_data[2602]=8'b01001111;
   assign rom_data[2603]=8'b10001001;
   assign rom_data[2604]=8'b01001111;
   assign rom_data[2605]=8'b10001001;
   assign rom_data[2606]=8'b01001111;
   assign rom_data[2607]=8'b10001001;
   assign rom_data[2608]=8'b01001111;
   assign rom_data[2609]=8'b10001010;
   assign rom_data[2610]=8'b01001111;
   assign rom_data[2611]=8'b10001010;
   assign rom_data[2612]=8'b01001111;
   assign rom_data[2613]=8'b10001010;
   assign rom_data[2614]=8'b01001111;
   assign rom_data[2615]=8'b10001010;
   assign rom_data[2616]=8'b01001111;
   assign rom_data[2617]=8'b10001010;
   assign rom_data[2618]=8'b01001111;
   assign rom_data[2619]=8'b10001001;
   assign rom_data[2620]=8'b01001111;
   assign rom_data[2621]=8'b10001001;
   assign rom_data[2622]=8'b01001111;
   assign rom_data[2623]=8'b10001001;
   assign rom_data[2624]=8'b01001111;
   assign rom_data[2625]=8'b10001000;
   assign rom_data[2626]=8'b01001111;
   assign rom_data[2627]=8'b10001000;
   assign rom_data[2628]=8'b01001111;
   assign rom_data[2629]=8'b10000111;
   assign rom_data[2630]=8'b01001111;
   assign rom_data[2631]=8'b10000111;
   assign rom_data[2632]=8'b01001111;
   assign rom_data[2633]=8'b10000110;
   assign rom_data[2634]=8'b01001111;
   assign rom_data[2635]=8'b10000101;
   assign rom_data[2636]=8'b01001111;
   assign rom_data[2637]=8'b10000100;
   assign rom_data[2638]=8'b01001111;
   assign rom_data[2639]=8'b10000011;
   assign rom_data[2640]=8'b01001111;
   assign rom_data[2641]=8'b10000011;
   assign rom_data[2642]=8'b01001111;
   assign rom_data[2643]=8'b10000010;
   assign rom_data[2644]=8'b01001111;
   assign rom_data[2645]=8'b10000001;
   assign rom_data[2646]=8'b01001111;
   assign rom_data[2647]=8'b10000000;
   assign rom_data[2648]=8'b01001111;
   assign rom_data[2649]=8'b01111110;
   assign rom_data[2650]=8'b01001111;
   assign rom_data[2651]=8'b01111101;
   assign rom_data[2652]=8'b01001111;
   assign rom_data[2653]=8'b01111100;
   assign rom_data[2654]=8'b01010000;
   assign rom_data[2655]=8'b01111011;
   assign rom_data[2656]=8'b01010000;
   assign rom_data[2657]=8'b01111010;
   assign rom_data[2658]=8'b01010000;
   assign rom_data[2659]=8'b01111001;
   assign rom_data[2660]=8'b01010000;
   assign rom_data[2661]=8'b01110111;
   assign rom_data[2662]=8'b01010000;
   assign rom_data[2663]=8'b01110110;
   assign rom_data[2664]=8'b01010000;
   assign rom_data[2665]=8'b01110101;
   assign rom_data[2666]=8'b01010000;
   assign rom_data[2667]=8'b01110100;
   assign rom_data[2668]=8'b01010000;
   assign rom_data[2669]=8'b01110010;
   assign rom_data[2670]=8'b01010000;
   assign rom_data[2671]=8'b01110001;
   assign rom_data[2672]=8'b01010000;
   assign rom_data[2673]=8'b01110000;
   assign rom_data[2674]=8'b01010000;
   assign rom_data[2675]=8'b01101110;
   assign rom_data[2676]=8'b01010000;
   assign rom_data[2677]=8'b01101101;
   assign rom_data[2678]=8'b01010000;
   assign rom_data[2679]=8'b01101100;
   assign rom_data[2680]=8'b01010000;
   assign rom_data[2681]=8'b01101010;
   assign rom_data[2682]=8'b01010000;
   assign rom_data[2683]=8'b01101001;
   assign rom_data[2684]=8'b01010000;
   assign rom_data[2685]=8'b01100111;
   assign rom_data[2686]=8'b01010000;
   assign rom_data[2687]=8'b01100110;
   assign rom_data[2688]=8'b01010000;
   assign rom_data[2689]=8'b01100101;
   assign rom_data[2690]=8'b01010000;
   assign rom_data[2691]=8'b01100011;
   assign rom_data[2692]=8'b01010000;
   assign rom_data[2693]=8'b01100010;
   assign rom_data[2694]=8'b01010000;
   assign rom_data[2695]=8'b01100001;
   assign rom_data[2696]=8'b01010000;
   assign rom_data[2697]=8'b01011111;
   assign rom_data[2698]=8'b01010000;
   assign rom_data[2699]=8'b01011110;
   assign rom_data[2700]=8'b01010000;
   assign rom_data[2701]=8'b01011100;
   assign rom_data[2702]=8'b01010000;
   assign rom_data[2703]=8'b01011011;
   assign rom_data[2704]=8'b01010000;
   assign rom_data[2705]=8'b01011001;
   assign rom_data[2706]=8'b01010000;
   assign rom_data[2707]=8'b01011000;
   assign rom_data[2708]=8'b01010000;
   assign rom_data[2709]=8'b01010111;
   assign rom_data[2710]=8'b01010000;
   assign rom_data[2711]=8'b01010101;
   assign rom_data[2712]=8'b01010000;
   assign rom_data[2713]=8'b01010100;
   assign rom_data[2714]=8'b01010000;
   assign rom_data[2715]=8'b01010010;
   assign rom_data[2716]=8'b01010000;
   assign rom_data[2717]=8'b01010001;
   assign rom_data[2718]=8'b01010000;
   assign rom_data[2719]=8'b01010000;
   assign rom_data[2720]=8'b01010000;
   assign rom_data[2721]=8'b01001110;
   assign rom_data[2722]=8'b01010000;
   assign rom_data[2723]=8'b01001101;
   assign rom_data[2724]=8'b01010000;
   assign rom_data[2725]=8'b01001100;
   assign rom_data[2726]=8'b01010000;
   assign rom_data[2727]=8'b01001010;
   assign rom_data[2728]=8'b01010000;
   assign rom_data[2729]=8'b01001001;
   assign rom_data[2730]=8'b01010000;
   assign rom_data[2731]=8'b01001000;
   assign rom_data[2732]=8'b01010000;
   assign rom_data[2733]=8'b01000110;
   assign rom_data[2734]=8'b01010000;
   assign rom_data[2735]=8'b01000101;
   assign rom_data[2736]=8'b01010000;
   assign rom_data[2737]=8'b01000100;
   assign rom_data[2738]=8'b01010001;
   assign rom_data[2739]=8'b01000010;
   assign rom_data[2740]=8'b01010001;
   assign rom_data[2741]=8'b01000001;
   assign rom_data[2742]=8'b01010001;
   assign rom_data[2743]=8'b01000000;
   assign rom_data[2744]=8'b01010001;
   assign rom_data[2745]=8'b00111111;
   assign rom_data[2746]=8'b01010001;
   assign rom_data[2747]=8'b00111101;
   assign rom_data[2748]=8'b01010001;
   assign rom_data[2749]=8'b00111100;
   assign rom_data[2750]=8'b01010001;
   assign rom_data[2751]=8'b00111011;
   assign rom_data[2752]=8'b01010001;
   assign rom_data[2753]=8'b00111010;
   assign rom_data[2754]=8'b01010001;
   assign rom_data[2755]=8'b00111001;
   assign rom_data[2756]=8'b01010001;
   assign rom_data[2757]=8'b00111000;
   assign rom_data[2758]=8'b01010001;
   assign rom_data[2759]=8'b00110110;
   assign rom_data[2760]=8'b01010001;
   assign rom_data[2761]=8'b00110101;
   assign rom_data[2762]=8'b01010001;
   assign rom_data[2763]=8'b00110100;
   assign rom_data[2764]=8'b01010001;
   assign rom_data[2765]=8'b00110011;
   assign rom_data[2766]=8'b01010001;
   assign rom_data[2767]=8'b00110011;
   assign rom_data[2768]=8'b01010001;
   assign rom_data[2769]=8'b00110010;
   assign rom_data[2770]=8'b01010001;
   assign rom_data[2771]=8'b00110001;
   assign rom_data[2772]=8'b01010001;
   assign rom_data[2773]=8'b00110000;
   assign rom_data[2774]=8'b01010001;
   assign rom_data[2775]=8'b00101111;
   assign rom_data[2776]=8'b01010001;
   assign rom_data[2777]=8'b00101111;
   assign rom_data[2778]=8'b01010001;
   assign rom_data[2779]=8'b00101110;
   assign rom_data[2780]=8'b01010001;
   assign rom_data[2781]=8'b00101110;
   assign rom_data[2782]=8'b01010001;
   assign rom_data[2783]=8'b00101101;
   assign rom_data[2784]=8'b01010001;
   assign rom_data[2785]=8'b00101101;
   assign rom_data[2786]=8'b01010001;
   assign rom_data[2787]=8'b00101100;
   assign rom_data[2788]=8'b01010001;
   assign rom_data[2789]=8'b00101100;
   assign rom_data[2790]=8'b01010001;
   assign rom_data[2791]=8'b00101100;
   assign rom_data[2792]=8'b01010001;
   assign rom_data[2793]=8'b00101100;
   assign rom_data[2794]=8'b01010001;
   assign rom_data[2795]=8'b00101100;
   assign rom_data[2796]=8'b01010001;
   assign rom_data[2797]=8'b00101100;
   assign rom_data[2798]=8'b01010001;
   assign rom_data[2799]=8'b00101100;
   assign rom_data[2800]=8'b01010001;
   assign rom_data[2801]=8'b00101101;
   assign rom_data[2802]=8'b01010001;
   assign rom_data[2803]=8'b00101101;
   assign rom_data[2804]=8'b01010001;
   assign rom_data[2805]=8'b00101101;
   assign rom_data[2806]=8'b01010010;
   assign rom_data[2807]=8'b00101110;
   assign rom_data[2808]=8'b01010010;
   assign rom_data[2809]=8'b00101111;
   assign rom_data[2810]=8'b01010010;
   assign rom_data[2811]=8'b00101111;
   assign rom_data[2812]=8'b01010010;
   assign rom_data[2813]=8'b00110000;
   assign rom_data[2814]=8'b01010010;
   assign rom_data[2815]=8'b00110001;
   assign rom_data[2816]=8'b01010010;
   assign rom_data[2817]=8'b00110001;
   assign rom_data[2818]=8'b01010010;
   assign rom_data[2819]=8'b00110010;
   assign rom_data[2820]=8'b01010010;
   assign rom_data[2821]=8'b00110011;
   assign rom_data[2822]=8'b01010010;
   assign rom_data[2823]=8'b00110100;
   assign rom_data[2824]=8'b01010010;
   assign rom_data[2825]=8'b00110101;
   assign rom_data[2826]=8'b01010010;
   assign rom_data[2827]=8'b00110110;
   assign rom_data[2828]=8'b01010010;
   assign rom_data[2829]=8'b00110111;
   assign rom_data[2830]=8'b01010010;
   assign rom_data[2831]=8'b00111000;
   assign rom_data[2832]=8'b01010010;
   assign rom_data[2833]=8'b00111010;
   assign rom_data[2834]=8'b01010010;
   assign rom_data[2835]=8'b00111011;
   assign rom_data[2836]=8'b01010010;
   assign rom_data[2837]=8'b00111100;
   assign rom_data[2838]=8'b01010010;
   assign rom_data[2839]=8'b00111101;
   assign rom_data[2840]=8'b01010010;
   assign rom_data[2841]=8'b00111110;
   assign rom_data[2842]=8'b01010010;
   assign rom_data[2843]=8'b01000000;
   assign rom_data[2844]=8'b01010010;
   assign rom_data[2845]=8'b01000001;
   assign rom_data[2846]=8'b01010010;
   assign rom_data[2847]=8'b01000010;
   assign rom_data[2848]=8'b01010010;
   assign rom_data[2849]=8'b01000100;
   assign rom_data[2850]=8'b01010010;
   assign rom_data[2851]=8'b01000101;
   assign rom_data[2852]=8'b01010010;
   assign rom_data[2853]=8'b01000110;
   assign rom_data[2854]=8'b01010010;
   assign rom_data[2855]=8'b01000111;
   assign rom_data[2856]=8'b01010010;
   assign rom_data[2857]=8'b01001001;
   assign rom_data[2858]=8'b01010010;
   assign rom_data[2859]=8'b01001010;
   assign rom_data[2860]=8'b01010010;
   assign rom_data[2861]=8'b01001100;
   assign rom_data[2862]=8'b01010010;
   assign rom_data[2863]=8'b01001101;
   assign rom_data[2864]=8'b01010010;
   assign rom_data[2865]=8'b01001110;
   assign rom_data[2866]=8'b01010010;
   assign rom_data[2867]=8'b01010000;
   assign rom_data[2868]=8'b01010010;
   assign rom_data[2869]=8'b01010001;
   assign rom_data[2870]=8'b01010010;
   assign rom_data[2871]=8'b01010010;
   assign rom_data[2872]=8'b01010010;
   assign rom_data[2873]=8'b01010100;
   assign rom_data[2874]=8'b01010010;
   assign rom_data[2875]=8'b01010101;
   assign rom_data[2876]=8'b01010010;
   assign rom_data[2877]=8'b01010111;
   assign rom_data[2878]=8'b01010010;
   assign rom_data[2879]=8'b01011000;
   assign rom_data[2880]=8'b01010010;
   assign rom_data[2881]=8'b01011010;
   assign rom_data[2882]=8'b01010011;
   assign rom_data[2883]=8'b01011011;
   assign rom_data[2884]=8'b01010011;
   assign rom_data[2885]=8'b01011100;
   assign rom_data[2886]=8'b01010011;
   assign rom_data[2887]=8'b01011110;
   assign rom_data[2888]=8'b01010011;
   assign rom_data[2889]=8'b01011111;
   assign rom_data[2890]=8'b01010011;
   assign rom_data[2891]=8'b01100001;
   assign rom_data[2892]=8'b01010011;
   assign rom_data[2893]=8'b01100010;
   assign rom_data[2894]=8'b01010011;
   assign rom_data[2895]=8'b01100011;
   assign rom_data[2896]=8'b01010011;
   assign rom_data[2897]=8'b01100101;
   assign rom_data[2898]=8'b01010011;
   assign rom_data[2899]=8'b01100110;
   assign rom_data[2900]=8'b01010011;
   assign rom_data[2901]=8'b01100111;
   assign rom_data[2902]=8'b01010011;
   assign rom_data[2903]=8'b01101001;
   assign rom_data[2904]=8'b01010011;
   assign rom_data[2905]=8'b01101010;
   assign rom_data[2906]=8'b01010011;
   assign rom_data[2907]=8'b01101100;
   assign rom_data[2908]=8'b01010011;
   assign rom_data[2909]=8'b01101101;
   assign rom_data[2910]=8'b01010011;
   assign rom_data[2911]=8'b01101110;
   assign rom_data[2912]=8'b01010011;
   assign rom_data[2913]=8'b01110000;
   assign rom_data[2914]=8'b01010011;
   assign rom_data[2915]=8'b01110001;
   assign rom_data[2916]=8'b01010011;
   assign rom_data[2917]=8'b01110010;
   assign rom_data[2918]=8'b01010011;
   assign rom_data[2919]=8'b01110100;
   assign rom_data[2920]=8'b01010011;
   assign rom_data[2921]=8'b01110101;
   assign rom_data[2922]=8'b01010011;
   assign rom_data[2923]=8'b01110110;
   assign rom_data[2924]=8'b01010011;
   assign rom_data[2925]=8'b01110111;
   assign rom_data[2926]=8'b01010011;
   assign rom_data[2927]=8'b01111001;
   assign rom_data[2928]=8'b01010011;
   assign rom_data[2929]=8'b01111010;
   assign rom_data[2930]=8'b01010011;
   assign rom_data[2931]=8'b01111011;
   assign rom_data[2932]=8'b01010011;
   assign rom_data[2933]=8'b01111100;
   assign rom_data[2934]=8'b01010011;
   assign rom_data[2935]=8'b01111101;
   assign rom_data[2936]=8'b01010011;
   assign rom_data[2937]=8'b01111110;
   assign rom_data[2938]=8'b01010011;
   assign rom_data[2939]=8'b01111111;
   assign rom_data[2940]=8'b01010011;
   assign rom_data[2941]=8'b10000000;
   assign rom_data[2942]=8'b01010011;
   assign rom_data[2943]=8'b10000001;
   assign rom_data[2944]=8'b01010011;
   assign rom_data[2945]=8'b10000010;
   assign rom_data[2946]=8'b01010011;
   assign rom_data[2947]=8'b10000011;
   assign rom_data[2948]=8'b01010011;
   assign rom_data[2949]=8'b10000100;
   assign rom_data[2950]=8'b01010011;
   assign rom_data[2951]=8'b10000101;
   assign rom_data[2952]=8'b01010011;
   assign rom_data[2953]=8'b10000110;
   assign rom_data[2954]=8'b01010011;
   assign rom_data[2955]=8'b10000110;
   assign rom_data[2956]=8'b01010011;
   assign rom_data[2957]=8'b10000111;
   assign rom_data[2958]=8'b01010011;
   assign rom_data[2959]=8'b10001000;
   assign rom_data[2960]=8'b01010100;
   assign rom_data[2961]=8'b10001000;
   assign rom_data[2962]=8'b01010100;
   assign rom_data[2963]=8'b10001001;
   assign rom_data[2964]=8'b01010100;
   assign rom_data[2965]=8'b10001001;
   assign rom_data[2966]=8'b01010100;
   assign rom_data[2967]=8'b10001001;
   assign rom_data[2968]=8'b01010100;
   assign rom_data[2969]=8'b10001010;
   assign rom_data[2970]=8'b01010100;
   assign rom_data[2971]=8'b10001010;
   assign rom_data[2972]=8'b01010100;
   assign rom_data[2973]=8'b10001010;
   assign rom_data[2974]=8'b01010100;
   assign rom_data[2975]=8'b10001010;
   assign rom_data[2976]=8'b01010100;
   assign rom_data[2977]=8'b10001010;
   assign rom_data[2978]=8'b01010100;
   assign rom_data[2979]=8'b10001001;
   assign rom_data[2980]=8'b01010100;
   assign rom_data[2981]=8'b10001001;
   assign rom_data[2982]=8'b01010100;
   assign rom_data[2983]=8'b10001001;
   assign rom_data[2984]=8'b01010100;
   assign rom_data[2985]=8'b10001000;
   assign rom_data[2986]=8'b01010100;
   assign rom_data[2987]=8'b10001000;
   assign rom_data[2988]=8'b01010100;
   assign rom_data[2989]=8'b10000111;
   assign rom_data[2990]=8'b01010100;
   assign rom_data[2991]=8'b10000111;
   assign rom_data[2992]=8'b01010100;
   assign rom_data[2993]=8'b10000110;
   assign rom_data[2994]=8'b01010100;
   assign rom_data[2995]=8'b10000101;
   assign rom_data[2996]=8'b01010100;
   assign rom_data[2997]=8'b10000100;
   assign rom_data[2998]=8'b01010100;
   assign rom_data[2999]=8'b10000011;
   assign rom_data[3000]=8'b01010100;
   assign rom_data[3001]=8'b10000011;
   assign rom_data[3002]=8'b01010100;
   assign rom_data[3003]=8'b10000010;
   assign rom_data[3004]=8'b01010100;
   assign rom_data[3005]=8'b10000001;
   assign rom_data[3006]=8'b01010100;
   assign rom_data[3007]=8'b10000000;
   assign rom_data[3008]=8'b01010100;
   assign rom_data[3009]=8'b01111110;
   assign rom_data[3010]=8'b01010100;
   assign rom_data[3011]=8'b01111101;
   assign rom_data[3012]=8'b01010100;
   assign rom_data[3013]=8'b01111100;
   assign rom_data[3014]=8'b01010100;
   assign rom_data[3015]=8'b01111011;
   assign rom_data[3016]=8'b01010100;
   assign rom_data[3017]=8'b01111010;
   assign rom_data[3018]=8'b01010100;
   assign rom_data[3019]=8'b01111001;
   assign rom_data[3020]=8'b01010100;
   assign rom_data[3021]=8'b01110111;
   assign rom_data[3022]=8'b01010100;
   assign rom_data[3023]=8'b01110110;
   assign rom_data[3024]=8'b01010100;
   assign rom_data[3025]=8'b01110101;
   assign rom_data[3026]=8'b01010100;
   assign rom_data[3027]=8'b01110100;
   assign rom_data[3028]=8'b01010101;
   assign rom_data[3029]=8'b01110010;
   assign rom_data[3030]=8'b01010101;
   assign rom_data[3031]=8'b01110001;
   assign rom_data[3032]=8'b01010101;
   assign rom_data[3033]=8'b01110000;
   assign rom_data[3034]=8'b01010101;
   assign rom_data[3035]=8'b01101110;
   assign rom_data[3036]=8'b01010101;
   assign rom_data[3037]=8'b01101101;
   assign rom_data[3038]=8'b01010101;
   assign rom_data[3039]=8'b01101100;
   assign rom_data[3040]=8'b01010101;
   assign rom_data[3041]=8'b01101010;
   assign rom_data[3042]=8'b01010101;
   assign rom_data[3043]=8'b01101001;
   assign rom_data[3044]=8'b01010101;
   assign rom_data[3045]=8'b01100111;
   assign rom_data[3046]=8'b01010101;
   assign rom_data[3047]=8'b01100110;
   assign rom_data[3048]=8'b01010101;
   assign rom_data[3049]=8'b01100101;
   assign rom_data[3050]=8'b01010101;
   assign rom_data[3051]=8'b01100011;
   assign rom_data[3052]=8'b01010101;
   assign rom_data[3053]=8'b01100010;
   assign rom_data[3054]=8'b01010101;
   assign rom_data[3055]=8'b01100001;
   assign rom_data[3056]=8'b01010101;
   assign rom_data[3057]=8'b01011111;
   assign rom_data[3058]=8'b01010101;
   assign rom_data[3059]=8'b01011110;
   assign rom_data[3060]=8'b01010101;
   assign rom_data[3061]=8'b01011100;
   assign rom_data[3062]=8'b01010101;
   assign rom_data[3063]=8'b01011011;
   assign rom_data[3064]=8'b01010101;
   assign rom_data[3065]=8'b01011001;
   assign rom_data[3066]=8'b01010101;
   assign rom_data[3067]=8'b01011000;
   assign rom_data[3068]=8'b01010101;
   assign rom_data[3069]=8'b01010111;
   assign rom_data[3070]=8'b01010101;
   assign rom_data[3071]=8'b01010101;
   assign rom_data[3072]=8'b01010101;
   assign rom_data[3073]=8'b01010100;
   assign rom_data[3074]=8'b01010101;
   assign rom_data[3075]=8'b01010010;
   assign rom_data[3076]=8'b01010101;
   assign rom_data[3077]=8'b01010001;
   assign rom_data[3078]=8'b01010101;
   assign rom_data[3079]=8'b01010000;
   assign rom_data[3080]=8'b01010101;
   assign rom_data[3081]=8'b01001110;
   assign rom_data[3082]=8'b01010101;
   assign rom_data[3083]=8'b01001101;
   assign rom_data[3084]=8'b01010101;
   assign rom_data[3085]=8'b01001100;
   assign rom_data[3086]=8'b01010101;
   assign rom_data[3087]=8'b01001010;
   assign rom_data[3088]=8'b01010101;
   assign rom_data[3089]=8'b01001001;
   assign rom_data[3090]=8'b01010101;
   assign rom_data[3091]=8'b01001000;
   assign rom_data[3092]=8'b01010101;
   assign rom_data[3093]=8'b01000110;
   assign rom_data[3094]=8'b01010101;
   assign rom_data[3095]=8'b01000101;
   assign rom_data[3096]=8'b01010101;
   assign rom_data[3097]=8'b01000100;
   assign rom_data[3098]=8'b01010101;
   assign rom_data[3099]=8'b01000010;
   assign rom_data[3100]=8'b01010101;
   assign rom_data[3101]=8'b01000001;
   assign rom_data[3102]=8'b01010101;
   assign rom_data[3103]=8'b01000000;
   assign rom_data[3104]=8'b01010101;
   assign rom_data[3105]=8'b00111111;
   assign rom_data[3106]=8'b01010101;
   assign rom_data[3107]=8'b00111101;
   assign rom_data[3108]=8'b01010101;
   assign rom_data[3109]=8'b00111100;
   assign rom_data[3110]=8'b01010101;
   assign rom_data[3111]=8'b00111011;
   assign rom_data[3112]=8'b01010110;
   assign rom_data[3113]=8'b00111010;
   assign rom_data[3114]=8'b01010110;
   assign rom_data[3115]=8'b00111001;
   assign rom_data[3116]=8'b01010110;
   assign rom_data[3117]=8'b00111000;
   assign rom_data[3118]=8'b01010110;
   assign rom_data[3119]=8'b00110110;
   assign rom_data[3120]=8'b01010110;
   assign rom_data[3121]=8'b00110101;
   assign rom_data[3122]=8'b01010110;
   assign rom_data[3123]=8'b00110100;
   assign rom_data[3124]=8'b01010110;
   assign rom_data[3125]=8'b00110011;
   assign rom_data[3126]=8'b01010110;
   assign rom_data[3127]=8'b00110011;
   assign rom_data[3128]=8'b01010110;
   assign rom_data[3129]=8'b00110010;
   assign rom_data[3130]=8'b01010110;
   assign rom_data[3131]=8'b00110001;
   assign rom_data[3132]=8'b01010110;
   assign rom_data[3133]=8'b00110000;
   assign rom_data[3134]=8'b01010110;
   assign rom_data[3135]=8'b00101111;
   assign rom_data[3136]=8'b01010110;
   assign rom_data[3137]=8'b00101111;
   assign rom_data[3138]=8'b01010110;
   assign rom_data[3139]=8'b00101110;
   assign rom_data[3140]=8'b01010110;
   assign rom_data[3141]=8'b00101110;
   assign rom_data[3142]=8'b01010110;
   assign rom_data[3143]=8'b00101101;
   assign rom_data[3144]=8'b01010110;
   assign rom_data[3145]=8'b00101101;
   assign rom_data[3146]=8'b01010110;
   assign rom_data[3147]=8'b00101100;
   assign rom_data[3148]=8'b01010110;
   assign rom_data[3149]=8'b00101100;
   assign rom_data[3150]=8'b01010110;
   assign rom_data[3151]=8'b00101100;
   assign rom_data[3152]=8'b01010110;
   assign rom_data[3153]=8'b00101100;
   assign rom_data[3154]=8'b01010110;
   assign rom_data[3155]=8'b00101100;
   assign rom_data[3156]=8'b01010110;
   assign rom_data[3157]=8'b00101100;
   assign rom_data[3158]=8'b01010110;
   assign rom_data[3159]=8'b00101100;
   assign rom_data[3160]=8'b01010110;
   assign rom_data[3161]=8'b00101101;
   assign rom_data[3162]=8'b01010110;
   assign rom_data[3163]=8'b00101101;
   assign rom_data[3164]=8'b01010110;
   assign rom_data[3165]=8'b00101101;
   assign rom_data[3166]=8'b01010110;
   assign rom_data[3167]=8'b00101110;
   assign rom_data[3168]=8'b01010110;
   assign rom_data[3169]=8'b00101111;
   assign rom_data[3170]=8'b01010110;
   assign rom_data[3171]=8'b00101111;
   assign rom_data[3172]=8'b01010110;
   assign rom_data[3173]=8'b00110000;
   assign rom_data[3174]=8'b01010110;
   assign rom_data[3175]=8'b00110001;
   assign rom_data[3176]=8'b01010110;
   assign rom_data[3177]=8'b00110001;
   assign rom_data[3178]=8'b01010111;
   assign rom_data[3179]=8'b00110010;
   assign rom_data[3180]=8'b01010111;
   assign rom_data[3181]=8'b00110011;
   assign rom_data[3182]=8'b01010111;
   assign rom_data[3183]=8'b00110100;
   assign rom_data[3184]=8'b01010111;
   assign rom_data[3185]=8'b00110101;
   assign rom_data[3186]=8'b01010111;
   assign rom_data[3187]=8'b00110110;
   assign rom_data[3188]=8'b01010111;
   assign rom_data[3189]=8'b00110111;
   assign rom_data[3190]=8'b01010111;
   assign rom_data[3191]=8'b00111000;
   assign rom_data[3192]=8'b01010111;
   assign rom_data[3193]=8'b00111010;
   assign rom_data[3194]=8'b01010111;
   assign rom_data[3195]=8'b00111011;
   assign rom_data[3196]=8'b01010111;
   assign rom_data[3197]=8'b00111100;
   assign rom_data[3198]=8'b01010111;
   assign rom_data[3199]=8'b00111101;
   assign rom_data[3200]=8'b01010111;
   assign rom_data[3201]=8'b00111110;
   assign rom_data[3202]=8'b01010111;
   assign rom_data[3203]=8'b01000000;
   assign rom_data[3204]=8'b01010111;
   assign rom_data[3205]=8'b01000001;
   assign rom_data[3206]=8'b01010111;
   assign rom_data[3207]=8'b01000010;
   assign rom_data[3208]=8'b01010111;
   assign rom_data[3209]=8'b01000100;
   assign rom_data[3210]=8'b01010111;
   assign rom_data[3211]=8'b01000101;
   assign rom_data[3212]=8'b01010111;
   assign rom_data[3213]=8'b01000110;
   assign rom_data[3214]=8'b01010111;
   assign rom_data[3215]=8'b01001000;
   assign rom_data[3216]=8'b01010111;
   assign rom_data[3217]=8'b01001001;
   assign rom_data[3218]=8'b01010111;
   assign rom_data[3219]=8'b01001010;
   assign rom_data[3220]=8'b01010111;
   assign rom_data[3221]=8'b01001100;
   assign rom_data[3222]=8'b01010111;
   assign rom_data[3223]=8'b01001101;
   assign rom_data[3224]=8'b01010111;
   assign rom_data[3225]=8'b01001110;
   assign rom_data[3226]=8'b01010111;
   assign rom_data[3227]=8'b01010000;
   assign rom_data[3228]=8'b01010111;
   assign rom_data[3229]=8'b01010001;
   assign rom_data[3230]=8'b01010111;
   assign rom_data[3231]=8'b01010010;
   assign rom_data[3232]=8'b01010111;
   assign rom_data[3233]=8'b01010100;
   assign rom_data[3234]=8'b01010111;
   assign rom_data[3235]=8'b01010101;
   assign rom_data[3236]=8'b01010111;
   assign rom_data[3237]=8'b01010111;
   assign rom_data[3238]=8'b01010111;
   assign rom_data[3239]=8'b01011000;
   assign rom_data[3240]=8'b01010111;
   assign rom_data[3241]=8'b01011010;
   assign rom_data[3242]=8'b01010111;
   assign rom_data[3243]=8'b01011011;
   assign rom_data[3244]=8'b01010111;
   assign rom_data[3245]=8'b01011100;
   assign rom_data[3246]=8'b01010111;
   assign rom_data[3247]=8'b01011110;
   assign rom_data[3248]=8'b01010111;
   assign rom_data[3249]=8'b01011111;
   assign rom_data[3250]=8'b01010111;
   assign rom_data[3251]=8'b01100001;
   assign rom_data[3252]=8'b01010111;
   assign rom_data[3253]=8'b01100010;
   assign rom_data[3254]=8'b01010111;
   assign rom_data[3255]=8'b01100011;
   assign rom_data[3256]=8'b01010111;
   assign rom_data[3257]=8'b01100101;
   assign rom_data[3258]=8'b01010111;
   assign rom_data[3259]=8'b01100110;
   assign rom_data[3260]=8'b01011000;
   assign rom_data[3261]=8'b01100111;
   assign rom_data[3262]=8'b01011000;
   assign rom_data[3263]=8'b01101001;
   assign rom_data[3264]=8'b01011000;
   assign rom_data[3265]=8'b01101010;
   assign rom_data[3266]=8'b01011000;
   assign rom_data[3267]=8'b01101100;
   assign rom_data[3268]=8'b01011000;
   assign rom_data[3269]=8'b01101101;
   assign rom_data[3270]=8'b01011000;
   assign rom_data[3271]=8'b01101110;
   assign rom_data[3272]=8'b01011000;
   assign rom_data[3273]=8'b01110000;
   assign rom_data[3274]=8'b01011000;
   assign rom_data[3275]=8'b01110001;
   assign rom_data[3276]=8'b01011000;
   assign rom_data[3277]=8'b01110010;
   assign rom_data[3278]=8'b01011000;
   assign rom_data[3279]=8'b01110100;
   assign rom_data[3280]=8'b01011000;
   assign rom_data[3281]=8'b01110101;
   assign rom_data[3282]=8'b01011000;
   assign rom_data[3283]=8'b01110110;
   assign rom_data[3284]=8'b01011000;
   assign rom_data[3285]=8'b01110111;
   assign rom_data[3286]=8'b01011000;
   assign rom_data[3287]=8'b01111001;
   assign rom_data[3288]=8'b01011000;
   assign rom_data[3289]=8'b01111010;
   assign rom_data[3290]=8'b01011000;
   assign rom_data[3291]=8'b01111011;
   assign rom_data[3292]=8'b01011000;
   assign rom_data[3293]=8'b01111100;
   assign rom_data[3294]=8'b01011000;
   assign rom_data[3295]=8'b01111101;
   assign rom_data[3296]=8'b01011000;
   assign rom_data[3297]=8'b01111110;
   assign rom_data[3298]=8'b01011000;
   assign rom_data[3299]=8'b01111111;
   assign rom_data[3300]=8'b01011000;
   assign rom_data[3301]=8'b10000000;
   assign rom_data[3302]=8'b01011000;
   assign rom_data[3303]=8'b10000001;
   assign rom_data[3304]=8'b01011000;
   assign rom_data[3305]=8'b10000010;
   assign rom_data[3306]=8'b01011000;
   assign rom_data[3307]=8'b10000011;
   assign rom_data[3308]=8'b01011000;
   assign rom_data[3309]=8'b10000100;
   assign rom_data[3310]=8'b01011000;
   assign rom_data[3311]=8'b10000101;
   assign rom_data[3312]=8'b01011000;
   assign rom_data[3313]=8'b10000110;
   assign rom_data[3314]=8'b01011000;
   assign rom_data[3315]=8'b10000110;
   assign rom_data[3316]=8'b01011000;
   assign rom_data[3317]=8'b10000111;
   assign rom_data[3318]=8'b01011000;
   assign rom_data[3319]=8'b10001000;
   assign rom_data[3320]=8'b01011000;
   assign rom_data[3321]=8'b10001000;
   assign rom_data[3322]=8'b01011000;
   assign rom_data[3323]=8'b10001001;
   assign rom_data[3324]=8'b01011000;
   assign rom_data[3325]=8'b10001001;
   assign rom_data[3326]=8'b01011000;
   assign rom_data[3327]=8'b10001001;
   assign rom_data[3328]=8'b01011000;
   assign rom_data[3329]=8'b10001010;
   assign rom_data[3330]=8'b01011000;
   assign rom_data[3331]=8'b10001010;
   assign rom_data[3332]=8'b01011001;
   assign rom_data[3333]=8'b10001010;
   assign rom_data[3334]=8'b01011001;
   assign rom_data[3335]=8'b10001010;
   assign rom_data[3336]=8'b01011001;
   assign rom_data[3337]=8'b10001010;
   assign rom_data[3338]=8'b01011001;
   assign rom_data[3339]=8'b10001001;
   assign rom_data[3340]=8'b01011001;
   assign rom_data[3341]=8'b10001001;
   assign rom_data[3342]=8'b01011001;
   assign rom_data[3343]=8'b10001001;
   assign rom_data[3344]=8'b01011001;
   assign rom_data[3345]=8'b10001000;
   assign rom_data[3346]=8'b01011001;
   assign rom_data[3347]=8'b10001000;
   assign rom_data[3348]=8'b01011001;
   assign rom_data[3349]=8'b10000111;
   assign rom_data[3350]=8'b01011001;
   assign rom_data[3351]=8'b10000111;
   assign rom_data[3352]=8'b01011001;
   assign rom_data[3353]=8'b10000110;
   assign rom_data[3354]=8'b01011001;
   assign rom_data[3355]=8'b10000101;
   assign rom_data[3356]=8'b01011001;
   assign rom_data[3357]=8'b10000100;
   assign rom_data[3358]=8'b01011001;
   assign rom_data[3359]=8'b10000011;
   assign rom_data[3360]=8'b01011001;
   assign rom_data[3361]=8'b10000011;
   assign rom_data[3362]=8'b01011001;
   assign rom_data[3363]=8'b10000010;
   assign rom_data[3364]=8'b01011001;
   assign rom_data[3365]=8'b10000001;
   assign rom_data[3366]=8'b01011001;
   assign rom_data[3367]=8'b10000000;
   assign rom_data[3368]=8'b01011001;
   assign rom_data[3369]=8'b01111110;
   assign rom_data[3370]=8'b01011001;
   assign rom_data[3371]=8'b01111101;
   assign rom_data[3372]=8'b01011001;
   assign rom_data[3373]=8'b01111100;
   assign rom_data[3374]=8'b01011001;
   assign rom_data[3375]=8'b01111011;
   assign rom_data[3376]=8'b01011001;
   assign rom_data[3377]=8'b01111010;
   assign rom_data[3378]=8'b01011001;
   assign rom_data[3379]=8'b01111001;
   assign rom_data[3380]=8'b01011001;
   assign rom_data[3381]=8'b01110111;
   assign rom_data[3382]=8'b01011001;
   assign rom_data[3383]=8'b01110110;
   assign rom_data[3384]=8'b01011001;
   assign rom_data[3385]=8'b01110101;
   assign rom_data[3386]=8'b01011001;
   assign rom_data[3387]=8'b01110100;
   assign rom_data[3388]=8'b01011001;
   assign rom_data[3389]=8'b01110010;
   assign rom_data[3390]=8'b01011001;
   assign rom_data[3391]=8'b01110001;
   assign rom_data[3392]=8'b01011001;
   assign rom_data[3393]=8'b01110000;
   assign rom_data[3394]=8'b01011001;
   assign rom_data[3395]=8'b01101110;
   assign rom_data[3396]=8'b01011001;
   assign rom_data[3397]=8'b01101101;
   assign rom_data[3398]=8'b01011001;
   assign rom_data[3399]=8'b01101100;
   assign rom_data[3400]=8'b01011001;
   assign rom_data[3401]=8'b01101010;
   assign rom_data[3402]=8'b01011001;
   assign rom_data[3403]=8'b01101001;
   assign rom_data[3404]=8'b01011010;
   assign rom_data[3405]=8'b01100111;
   assign rom_data[3406]=8'b01011010;
   assign rom_data[3407]=8'b01100110;
   assign rom_data[3408]=8'b01011010;
   assign rom_data[3409]=8'b01100101;
   assign rom_data[3410]=8'b01011010;
   assign rom_data[3411]=8'b01100011;
   assign rom_data[3412]=8'b01011010;
   assign rom_data[3413]=8'b01100010;
   assign rom_data[3414]=8'b01011010;
   assign rom_data[3415]=8'b01100001;
   assign rom_data[3416]=8'b01011010;
   assign rom_data[3417]=8'b01011111;
   assign rom_data[3418]=8'b01011010;
   assign rom_data[3419]=8'b01011110;
   assign rom_data[3420]=8'b01011010;
   assign rom_data[3421]=8'b01011100;
   assign rom_data[3422]=8'b01011010;
   assign rom_data[3423]=8'b01011011;
   assign rom_data[3424]=8'b01011010;
   assign rom_data[3425]=8'b01011001;
   assign rom_data[3426]=8'b01011010;
   assign rom_data[3427]=8'b01011000;
   assign rom_data[3428]=8'b01011010;
   assign rom_data[3429]=8'b01010111;
   assign rom_data[3430]=8'b01011010;
   assign rom_data[3431]=8'b01010101;
   assign rom_data[3432]=8'b01011010;
   assign rom_data[3433]=8'b01010100;
   assign rom_data[3434]=8'b01011010;
   assign rom_data[3435]=8'b01010010;
   assign rom_data[3436]=8'b01011010;
   assign rom_data[3437]=8'b01010001;
   assign rom_data[3438]=8'b01011010;
   assign rom_data[3439]=8'b01010000;
   assign rom_data[3440]=8'b01011010;
   assign rom_data[3441]=8'b01001110;
   assign rom_data[3442]=8'b01011010;
   assign rom_data[3443]=8'b01001101;
   assign rom_data[3444]=8'b01011010;
   assign rom_data[3445]=8'b01001100;
   assign rom_data[3446]=8'b01011010;
   assign rom_data[3447]=8'b01001010;
   assign rom_data[3448]=8'b01011010;
   assign rom_data[3449]=8'b01001001;
   assign rom_data[3450]=8'b01011010;
   assign rom_data[3451]=8'b01001000;
   assign rom_data[3452]=8'b01011010;
   assign rom_data[3453]=8'b01000110;
   assign rom_data[3454]=8'b01011010;
   assign rom_data[3455]=8'b01000101;
   assign rom_data[3456]=8'b01011010;
   assign rom_data[3457]=8'b01000100;
   assign rom_data[3458]=8'b01011010;
   assign rom_data[3459]=8'b01000010;
   assign rom_data[3460]=8'b01011010;
   assign rom_data[3461]=8'b01000001;
   assign rom_data[3462]=8'b01011010;
   assign rom_data[3463]=8'b01000000;
   assign rom_data[3464]=8'b01011010;
   assign rom_data[3465]=8'b00111111;
   assign rom_data[3466]=8'b01011010;
   assign rom_data[3467]=8'b00111101;
   assign rom_data[3468]=8'b01011010;
   assign rom_data[3469]=8'b00111100;
   assign rom_data[3470]=8'b01011010;
   assign rom_data[3471]=8'b00111011;
   assign rom_data[3472]=8'b01011010;
   assign rom_data[3473]=8'b00111010;
   assign rom_data[3474]=8'b01011010;
   assign rom_data[3475]=8'b00111001;
   assign rom_data[3476]=8'b01011010;
   assign rom_data[3477]=8'b00111000;
   assign rom_data[3478]=8'b01011010;
   assign rom_data[3479]=8'b00110110;
   assign rom_data[3480]=8'b01011010;
   assign rom_data[3481]=8'b00110101;
   assign rom_data[3482]=8'b01011010;
   assign rom_data[3483]=8'b00110100;
   assign rom_data[3484]=8'b01011010;
   assign rom_data[3485]=8'b00110011;
   assign rom_data[3486]=8'b01011011;
   assign rom_data[3487]=8'b00110011;
   assign rom_data[3488]=8'b01011011;
   assign rom_data[3489]=8'b00110010;
   assign rom_data[3490]=8'b01011011;
   assign rom_data[3491]=8'b00110001;
   assign rom_data[3492]=8'b01011011;
   assign rom_data[3493]=8'b00110000;
   assign rom_data[3494]=8'b01011011;
   assign rom_data[3495]=8'b00101111;
   assign rom_data[3496]=8'b01011011;
   assign rom_data[3497]=8'b00101111;
   assign rom_data[3498]=8'b01011011;
   assign rom_data[3499]=8'b00101110;
   assign rom_data[3500]=8'b01011011;
   assign rom_data[3501]=8'b00101110;
   assign rom_data[3502]=8'b01011011;
   assign rom_data[3503]=8'b00101101;
   assign rom_data[3504]=8'b01011011;
   assign rom_data[3505]=8'b00101101;
   assign rom_data[3506]=8'b01011011;
   assign rom_data[3507]=8'b00101100;
   assign rom_data[3508]=8'b01011011;
   assign rom_data[3509]=8'b00101100;
   assign rom_data[3510]=8'b01011011;
   assign rom_data[3511]=8'b00101100;
   assign rom_data[3512]=8'b01011011;
   assign rom_data[3513]=8'b00101100;
   assign rom_data[3514]=8'b01011011;
   assign rom_data[3515]=8'b00101100;
   assign rom_data[3516]=8'b01011011;
   assign rom_data[3517]=8'b00101100;
   assign rom_data[3518]=8'b01011011;
   assign rom_data[3519]=8'b00101100;
   assign rom_data[3520]=8'b01011011;
   assign rom_data[3521]=8'b00101101;
   assign rom_data[3522]=8'b01011011;
   assign rom_data[3523]=8'b00101101;
   assign rom_data[3524]=8'b01011011;
   assign rom_data[3525]=8'b00101101;
   assign rom_data[3526]=8'b01011011;
   assign rom_data[3527]=8'b00101110;
   assign rom_data[3528]=8'b01011011;
   assign rom_data[3529]=8'b00101111;
   assign rom_data[3530]=8'b01011011;
   assign rom_data[3531]=8'b00101111;
   assign rom_data[3532]=8'b01011011;
   assign rom_data[3533]=8'b00110000;
   assign rom_data[3534]=8'b01011011;
   assign rom_data[3535]=8'b00110001;
   assign rom_data[3536]=8'b01011011;
   assign rom_data[3537]=8'b00110001;
   assign rom_data[3538]=8'b01011011;
   assign rom_data[3539]=8'b00110010;
   assign rom_data[3540]=8'b01011011;
   assign rom_data[3541]=8'b00110011;
   assign rom_data[3542]=8'b01011011;
   assign rom_data[3543]=8'b00110100;
   assign rom_data[3544]=8'b01011011;
   assign rom_data[3545]=8'b00110101;
   assign rom_data[3546]=8'b01011011;
   assign rom_data[3547]=8'b00110110;
   assign rom_data[3548]=8'b01011011;
   assign rom_data[3549]=8'b00110111;
   assign rom_data[3550]=8'b01011011;
   assign rom_data[3551]=8'b00111000;
   assign rom_data[3552]=8'b01011100;
   assign rom_data[3553]=8'b00111010;
   assign rom_data[3554]=8'b01011100;
   assign rom_data[3555]=8'b00111011;
   assign rom_data[3556]=8'b01011100;
   assign rom_data[3557]=8'b00111100;
   assign rom_data[3558]=8'b01011100;
   assign rom_data[3559]=8'b00111101;
   assign rom_data[3560]=8'b01011100;
   assign rom_data[3561]=8'b00111110;
   assign rom_data[3562]=8'b01011100;
   assign rom_data[3563]=8'b01000000;
   assign rom_data[3564]=8'b01011100;
   assign rom_data[3565]=8'b01000001;
   assign rom_data[3566]=8'b01011100;
   assign rom_data[3567]=8'b01000010;
   assign rom_data[3568]=8'b01011100;
   assign rom_data[3569]=8'b01000100;
   assign rom_data[3570]=8'b01011100;
   assign rom_data[3571]=8'b01000101;
   assign rom_data[3572]=8'b01011100;
   assign rom_data[3573]=8'b01000110;
   assign rom_data[3574]=8'b01011100;
   assign rom_data[3575]=8'b01001000;
   assign rom_data[3576]=8'b01011100;
   assign rom_data[3577]=8'b01001001;
   assign rom_data[3578]=8'b01011100;
   assign rom_data[3579]=8'b01001010;
   assign rom_data[3580]=8'b01011100;
   assign rom_data[3581]=8'b01001100;
   assign rom_data[3582]=8'b01011100;
   assign rom_data[3583]=8'b01001101;
   assign rom_data[3584]=8'b01011100;
   assign rom_data[3585]=8'b01001110;
   assign rom_data[3586]=8'b01011100;
   assign rom_data[3587]=8'b01010000;
   assign rom_data[3588]=8'b01011100;
   assign rom_data[3589]=8'b01010001;
   assign rom_data[3590]=8'b01011100;
   assign rom_data[3591]=8'b01010011;
   assign rom_data[3592]=8'b01011100;
   assign rom_data[3593]=8'b01010100;
   assign rom_data[3594]=8'b01011100;
   assign rom_data[3595]=8'b01010101;
   assign rom_data[3596]=8'b01011100;
   assign rom_data[3597]=8'b01010111;
   assign rom_data[3598]=8'b01011100;
   assign rom_data[3599]=8'b01011000;
   assign rom_data[3600]=8'b01011100;
   assign rom_data[3601]=8'b01011010;
   assign rom_data[3602]=8'b01011100;
   assign rom_data[3603]=8'b01011011;
   assign rom_data[3604]=8'b01011100;
   assign rom_data[3605]=8'b01011100;
   assign rom_data[3606]=8'b01011100;
   assign rom_data[3607]=8'b01011110;
   assign rom_data[3608]=8'b01011100;
   assign rom_data[3609]=8'b01011111;
   assign rom_data[3610]=8'b01011100;
   assign rom_data[3611]=8'b01100001;
   assign rom_data[3612]=8'b01011100;
   assign rom_data[3613]=8'b01100010;
   assign rom_data[3614]=8'b01011100;
   assign rom_data[3615]=8'b01100011;
   assign rom_data[3616]=8'b01011100;
   assign rom_data[3617]=8'b01100101;
   assign rom_data[3618]=8'b01011100;
   assign rom_data[3619]=8'b01100110;
   assign rom_data[3620]=8'b01011100;
   assign rom_data[3621]=8'b01100111;
   assign rom_data[3622]=8'b01011100;
   assign rom_data[3623]=8'b01101001;
   assign rom_data[3624]=8'b01011100;
   assign rom_data[3625]=8'b01101010;
   assign rom_data[3626]=8'b01011100;
   assign rom_data[3627]=8'b01101100;
   assign rom_data[3628]=8'b01011100;
   assign rom_data[3629]=8'b01101101;
   assign rom_data[3630]=8'b01011100;
   assign rom_data[3631]=8'b01101110;
   assign rom_data[3632]=8'b01011100;
   assign rom_data[3633]=8'b01110000;
   assign rom_data[3634]=8'b01011100;
   assign rom_data[3635]=8'b01110001;
   assign rom_data[3636]=8'b01011101;
   assign rom_data[3637]=8'b01110010;
   assign rom_data[3638]=8'b01011101;
   assign rom_data[3639]=8'b01110100;
   assign rom_data[3640]=8'b01011101;
   assign rom_data[3641]=8'b01110101;
   assign rom_data[3642]=8'b01011101;
   assign rom_data[3643]=8'b01110110;
   assign rom_data[3644]=8'b01011101;
   assign rom_data[3645]=8'b01110111;
   assign rom_data[3646]=8'b01011101;
   assign rom_data[3647]=8'b01111001;
   assign rom_data[3648]=8'b01011101;
   assign rom_data[3649]=8'b01111010;
   assign rom_data[3650]=8'b01011101;
   assign rom_data[3651]=8'b01111011;
   assign rom_data[3652]=8'b01011101;
   assign rom_data[3653]=8'b01111100;
   assign rom_data[3654]=8'b01011101;
   assign rom_data[3655]=8'b01111101;
   assign rom_data[3656]=8'b01011101;
   assign rom_data[3657]=8'b01111110;
   assign rom_data[3658]=8'b01011101;
   assign rom_data[3659]=8'b01111111;
   assign rom_data[3660]=8'b01011101;
   assign rom_data[3661]=8'b10000000;
   assign rom_data[3662]=8'b01011101;
   assign rom_data[3663]=8'b10000001;
   assign rom_data[3664]=8'b01011101;
   assign rom_data[3665]=8'b10000010;
   assign rom_data[3666]=8'b01011101;
   assign rom_data[3667]=8'b10000011;
   assign rom_data[3668]=8'b01011101;
   assign rom_data[3669]=8'b10000100;
   assign rom_data[3670]=8'b01011101;
   assign rom_data[3671]=8'b10000101;
   assign rom_data[3672]=8'b01011101;
   assign rom_data[3673]=8'b10000110;
   assign rom_data[3674]=8'b01011101;
   assign rom_data[3675]=8'b10000110;
   assign rom_data[3676]=8'b01011101;
   assign rom_data[3677]=8'b10000111;
   assign rom_data[3678]=8'b01011101;
   assign rom_data[3679]=8'b10001000;
   assign rom_data[3680]=8'b01011101;
   assign rom_data[3681]=8'b10001000;
   assign rom_data[3682]=8'b01011101;
   assign rom_data[3683]=8'b10001001;
   assign rom_data[3684]=8'b01011101;
   assign rom_data[3685]=8'b10001001;
   assign rom_data[3686]=8'b01011101;
   assign rom_data[3687]=8'b10001001;
   assign rom_data[3688]=8'b01011101;
   assign rom_data[3689]=8'b10001010;
   assign rom_data[3690]=8'b01011101;
   assign rom_data[3691]=8'b10001010;
   assign rom_data[3692]=8'b01011101;
   assign rom_data[3693]=8'b10001010;
   assign rom_data[3694]=8'b01011101;
   assign rom_data[3695]=8'b10001010;
   assign rom_data[3696]=8'b01011101;
   assign rom_data[3697]=8'b10001010;
   assign rom_data[3698]=8'b01011101;
   assign rom_data[3699]=8'b10001001;
   assign rom_data[3700]=8'b01011101;
   assign rom_data[3701]=8'b10001001;
   assign rom_data[3702]=8'b01011101;
   assign rom_data[3703]=8'b10001001;
   assign rom_data[3704]=8'b01011110;
   assign rom_data[3705]=8'b10001000;
   assign rom_data[3706]=8'b01011110;
   assign rom_data[3707]=8'b10001000;
   assign rom_data[3708]=8'b01011110;
   assign rom_data[3709]=8'b10000111;
   assign rom_data[3710]=8'b01011110;
   assign rom_data[3711]=8'b10000111;
   assign rom_data[3712]=8'b01011110;
   assign rom_data[3713]=8'b10000110;
   assign rom_data[3714]=8'b01011110;
   assign rom_data[3715]=8'b10000101;
   assign rom_data[3716]=8'b01011110;
   assign rom_data[3717]=8'b10000100;
   assign rom_data[3718]=8'b01011110;
   assign rom_data[3719]=8'b10000011;
   assign rom_data[3720]=8'b01011110;
   assign rom_data[3721]=8'b10000011;
   assign rom_data[3722]=8'b01011110;
   assign rom_data[3723]=8'b10000010;
   assign rom_data[3724]=8'b01011110;
   assign rom_data[3725]=8'b10000001;
   assign rom_data[3726]=8'b01011110;
   assign rom_data[3727]=8'b10000000;
   assign rom_data[3728]=8'b01011110;
   assign rom_data[3729]=8'b01111110;
   assign rom_data[3730]=8'b01011110;
   assign rom_data[3731]=8'b01111101;
   assign rom_data[3732]=8'b01011110;
   assign rom_data[3733]=8'b01111100;
   assign rom_data[3734]=8'b01011110;
   assign rom_data[3735]=8'b01111011;
   assign rom_data[3736]=8'b01011110;
   assign rom_data[3737]=8'b01111010;
   assign rom_data[3738]=8'b01011110;
   assign rom_data[3739]=8'b01111001;
   assign rom_data[3740]=8'b01011110;
   assign rom_data[3741]=8'b01110111;
   assign rom_data[3742]=8'b01011110;
   assign rom_data[3743]=8'b01110110;
   assign rom_data[3744]=8'b01011110;
   assign rom_data[3745]=8'b01110101;
   assign rom_data[3746]=8'b01011110;
   assign rom_data[3747]=8'b01110100;
   assign rom_data[3748]=8'b01011110;
   assign rom_data[3749]=8'b01110010;
   assign rom_data[3750]=8'b01011110;
   assign rom_data[3751]=8'b01110001;
   assign rom_data[3752]=8'b01011110;
   assign rom_data[3753]=8'b01110000;
   assign rom_data[3754]=8'b01011110;
   assign rom_data[3755]=8'b01101110;
   assign rom_data[3756]=8'b01011110;
   assign rom_data[3757]=8'b01101101;
   assign rom_data[3758]=8'b01011110;
   assign rom_data[3759]=8'b01101100;
   assign rom_data[3760]=8'b01011110;
   assign rom_data[3761]=8'b01101010;
   assign rom_data[3762]=8'b01011110;
   assign rom_data[3763]=8'b01101001;
   assign rom_data[3764]=8'b01011110;
   assign rom_data[3765]=8'b01100111;
   assign rom_data[3766]=8'b01011110;
   assign rom_data[3767]=8'b01100110;
   assign rom_data[3768]=8'b01011110;
   assign rom_data[3769]=8'b01100101;
   assign rom_data[3770]=8'b01011110;
   assign rom_data[3771]=8'b01100011;
   assign rom_data[3772]=8'b01011110;
   assign rom_data[3773]=8'b01100010;
   assign rom_data[3774]=8'b01011110;
   assign rom_data[3775]=8'b01100001;
   assign rom_data[3776]=8'b01011110;
   assign rom_data[3777]=8'b01011111;
   assign rom_data[3778]=8'b01011110;
   assign rom_data[3779]=8'b01011110;
   assign rom_data[3780]=8'b01011111;
   assign rom_data[3781]=8'b01011100;
   assign rom_data[3782]=8'b01011111;
   assign rom_data[3783]=8'b01011011;
   assign rom_data[3784]=8'b01011111;
   assign rom_data[3785]=8'b01011001;
   assign rom_data[3786]=8'b01011111;
   assign rom_data[3787]=8'b01011000;
   assign rom_data[3788]=8'b01011111;
   assign rom_data[3789]=8'b01010111;
   assign rom_data[3790]=8'b01011111;
   assign rom_data[3791]=8'b01010101;
   assign rom_data[3792]=8'b01011111;
   assign rom_data[3793]=8'b01010100;
   assign rom_data[3794]=8'b01011111;
   assign rom_data[3795]=8'b01010010;
   assign rom_data[3796]=8'b01011111;
   assign rom_data[3797]=8'b01010001;
   assign rom_data[3798]=8'b01011111;
   assign rom_data[3799]=8'b01010000;
   assign rom_data[3800]=8'b01011111;
   assign rom_data[3801]=8'b01001110;
   assign rom_data[3802]=8'b01011111;
   assign rom_data[3803]=8'b01001101;
   assign rom_data[3804]=8'b01011111;
   assign rom_data[3805]=8'b01001100;
   assign rom_data[3806]=8'b01011111;
   assign rom_data[3807]=8'b01001010;
   assign rom_data[3808]=8'b01011111;
   assign rom_data[3809]=8'b01001001;
   assign rom_data[3810]=8'b01011111;
   assign rom_data[3811]=8'b01001000;
   assign rom_data[3812]=8'b01011111;
   assign rom_data[3813]=8'b01000110;
   assign rom_data[3814]=8'b01011111;
   assign rom_data[3815]=8'b01000101;
   assign rom_data[3816]=8'b01011111;
   assign rom_data[3817]=8'b01000100;
   assign rom_data[3818]=8'b01011111;
   assign rom_data[3819]=8'b01000010;
   assign rom_data[3820]=8'b01011111;
   assign rom_data[3821]=8'b01000001;
   assign rom_data[3822]=8'b01011111;
   assign rom_data[3823]=8'b01000000;
   assign rom_data[3824]=8'b01011111;
   assign rom_data[3825]=8'b00111111;
   assign rom_data[3826]=8'b01011111;
   assign rom_data[3827]=8'b00111101;
   assign rom_data[3828]=8'b01011111;
   assign rom_data[3829]=8'b00111100;
   assign rom_data[3830]=8'b01011111;
   assign rom_data[3831]=8'b00111011;
   assign rom_data[3832]=8'b01011111;
   assign rom_data[3833]=8'b00111010;
   assign rom_data[3834]=8'b01011111;
   assign rom_data[3835]=8'b00111001;
   assign rom_data[3836]=8'b01011111;
   assign rom_data[3837]=8'b00111000;
   assign rom_data[3838]=8'b01011111;
   assign rom_data[3839]=8'b00110110;
   assign rom_data[3840]=8'b01011111;
   assign rom_data[3841]=8'b00110101;
   assign rom_data[3842]=8'b01011111;
   assign rom_data[3843]=8'b00110100;
   assign rom_data[3844]=8'b01011111;
   assign rom_data[3845]=8'b00110011;
   assign rom_data[3846]=8'b01011111;
   assign rom_data[3847]=8'b00110011;
   assign rom_data[3848]=8'b01011111;
   assign rom_data[3849]=8'b00110010;
   assign rom_data[3850]=8'b01011111;
   assign rom_data[3851]=8'b00110001;
   assign rom_data[3852]=8'b01011111;
   assign rom_data[3853]=8'b00110000;
   assign rom_data[3854]=8'b01011111;
   assign rom_data[3855]=8'b00101111;
   assign rom_data[3856]=8'b01011111;
   assign rom_data[3857]=8'b00101111;
   assign rom_data[3858]=8'b01011111;
   assign rom_data[3859]=8'b00101110;
   assign rom_data[3860]=8'b01100000;
   assign rom_data[3861]=8'b00101110;
   assign rom_data[3862]=8'b01100000;
   assign rom_data[3863]=8'b00101101;
   assign rom_data[3864]=8'b01100000;
   assign rom_data[3865]=8'b00101101;
   assign rom_data[3866]=8'b01100000;
   assign rom_data[3867]=8'b00101100;
   assign rom_data[3868]=8'b01100000;
   assign rom_data[3869]=8'b00101100;
   assign rom_data[3870]=8'b01100000;
   assign rom_data[3871]=8'b00101100;
   assign rom_data[3872]=8'b01100000;
   assign rom_data[3873]=8'b00101100;
   assign rom_data[3874]=8'b01100000;
   assign rom_data[3875]=8'b00101100;
   assign rom_data[3876]=8'b01100000;
   assign rom_data[3877]=8'b00101100;
   assign rom_data[3878]=8'b01100000;
   assign rom_data[3879]=8'b00101100;
   assign rom_data[3880]=8'b01100000;
   assign rom_data[3881]=8'b00101101;
   assign rom_data[3882]=8'b01100000;
   assign rom_data[3883]=8'b00101101;
   assign rom_data[3884]=8'b01100000;
   assign rom_data[3885]=8'b00101101;
   assign rom_data[3886]=8'b01100000;
   assign rom_data[3887]=8'b00101110;
   assign rom_data[3888]=8'b01100000;
   assign rom_data[3889]=8'b00101111;
   assign rom_data[3890]=8'b01100000;
   assign rom_data[3891]=8'b00101111;
   assign rom_data[3892]=8'b01100000;
   assign rom_data[3893]=8'b00110000;
   assign rom_data[3894]=8'b01100000;
   assign rom_data[3895]=8'b00110001;
   assign rom_data[3896]=8'b01100000;
   assign rom_data[3897]=8'b00110001;
   assign rom_data[3898]=8'b01100000;
   assign rom_data[3899]=8'b00110010;
   assign rom_data[3900]=8'b01100000;
   assign rom_data[3901]=8'b00110011;
   assign rom_data[3902]=8'b01100000;
   assign rom_data[3903]=8'b00110100;
   assign rom_data[3904]=8'b01100000;
   assign rom_data[3905]=8'b00110101;
   assign rom_data[3906]=8'b01100000;
   assign rom_data[3907]=8'b00110110;
   assign rom_data[3908]=8'b01100000;
   assign rom_data[3909]=8'b00110111;
   assign rom_data[3910]=8'b01100000;
   assign rom_data[3911]=8'b00111000;
   assign rom_data[3912]=8'b01100000;
   assign rom_data[3913]=8'b00111010;
   assign rom_data[3914]=8'b01100000;
   assign rom_data[3915]=8'b00111011;
   assign rom_data[3916]=8'b01100000;
   assign rom_data[3917]=8'b00111100;
   assign rom_data[3918]=8'b01100000;
   assign rom_data[3919]=8'b00111101;
   assign rom_data[3920]=8'b01100000;
   assign rom_data[3921]=8'b00111110;
   assign rom_data[3922]=8'b01100000;
   assign rom_data[3923]=8'b01000000;
   assign rom_data[3924]=8'b01100000;
   assign rom_data[3925]=8'b01000001;
   assign rom_data[3926]=8'b01100001;
   assign rom_data[3927]=8'b01000010;
   assign rom_data[3928]=8'b01100001;
   assign rom_data[3929]=8'b01000100;
   assign rom_data[3930]=8'b01100001;
   assign rom_data[3931]=8'b01000101;
   assign rom_data[3932]=8'b01100001;
   assign rom_data[3933]=8'b01000110;
   assign rom_data[3934]=8'b01100001;
   assign rom_data[3935]=8'b01001000;
   assign rom_data[3936]=8'b01100001;
   assign rom_data[3937]=8'b01001001;
   assign rom_data[3938]=8'b01100001;
   assign rom_data[3939]=8'b01001010;
   assign rom_data[3940]=8'b01100001;
   assign rom_data[3941]=8'b01001100;
   assign rom_data[3942]=8'b01100001;
   assign rom_data[3943]=8'b01001101;
   assign rom_data[3944]=8'b01100001;
   assign rom_data[3945]=8'b01001110;
   assign rom_data[3946]=8'b01100001;
   assign rom_data[3947]=8'b01010000;
   assign rom_data[3948]=8'b01100001;
   assign rom_data[3949]=8'b01010001;
   assign rom_data[3950]=8'b01100001;
   assign rom_data[3951]=8'b01010011;
   assign rom_data[3952]=8'b01100001;
   assign rom_data[3953]=8'b01010100;
   assign rom_data[3954]=8'b01100001;
   assign rom_data[3955]=8'b01010101;
   assign rom_data[3956]=8'b01100001;
   assign rom_data[3957]=8'b01010111;
   assign rom_data[3958]=8'b01100001;
   assign rom_data[3959]=8'b01011000;
   assign rom_data[3960]=8'b01100001;
   assign rom_data[3961]=8'b01011010;
   assign rom_data[3962]=8'b01100001;
   assign rom_data[3963]=8'b01011011;
   assign rom_data[3964]=8'b01100001;
   assign rom_data[3965]=8'b01011100;
   assign rom_data[3966]=8'b01100001;
   assign rom_data[3967]=8'b01011110;
   assign rom_data[3968]=8'b01100001;
   assign rom_data[3969]=8'b01011111;
   assign rom_data[3970]=8'b01100001;
   assign rom_data[3971]=8'b01100001;
   assign rom_data[3972]=8'b01100001;
   assign rom_data[3973]=8'b01100010;
   assign rom_data[3974]=8'b01100001;
   assign rom_data[3975]=8'b01100011;
   assign rom_data[3976]=8'b01100001;
   assign rom_data[3977]=8'b01100101;
   assign rom_data[3978]=8'b01100001;
   assign rom_data[3979]=8'b01100110;
   assign rom_data[3980]=8'b01100001;
   assign rom_data[3981]=8'b01100111;
   assign rom_data[3982]=8'b01100001;
   assign rom_data[3983]=8'b01101001;
   assign rom_data[3984]=8'b01100001;
   assign rom_data[3985]=8'b01101010;
   assign rom_data[3986]=8'b01100001;
   assign rom_data[3987]=8'b01101100;
   assign rom_data[3988]=8'b01100001;
   assign rom_data[3989]=8'b01101101;
   assign rom_data[3990]=8'b01100001;
   assign rom_data[3991]=8'b01101110;
   assign rom_data[3992]=8'b01100001;
   assign rom_data[3993]=8'b01110000;
   assign rom_data[3994]=8'b01100001;
   assign rom_data[3995]=8'b01110001;
   assign rom_data[3996]=8'b01100001;
   assign rom_data[3997]=8'b01110010;
   assign rom_data[3998]=8'b01100001;
   assign rom_data[3999]=8'b01110100;
   assign rom_data[4000]=8'b01100001;
   assign rom_data[4001]=8'b01110101;
   assign rom_data[4002]=8'b01100001;
   assign rom_data[4003]=8'b01110110;
   assign rom_data[4004]=8'b01100001;
   assign rom_data[4005]=8'b01110111;
   assign rom_data[4006]=8'b01100001;
   assign rom_data[4007]=8'b01111001;
   assign rom_data[4008]=8'b01100001;
   assign rom_data[4009]=8'b01111010;
   assign rom_data[4010]=8'b01100010;
   assign rom_data[4011]=8'b01111011;
   assign rom_data[4012]=8'b01100010;
   assign rom_data[4013]=8'b01111100;
   assign rom_data[4014]=8'b01100010;
   assign rom_data[4015]=8'b01111101;
   assign rom_data[4016]=8'b01100010;
   assign rom_data[4017]=8'b01111110;
   assign rom_data[4018]=8'b01100010;
   assign rom_data[4019]=8'b01111111;
   assign rom_data[4020]=8'b01100010;
   assign rom_data[4021]=8'b10000000;
   assign rom_data[4022]=8'b01100010;
   assign rom_data[4023]=8'b10000001;
   assign rom_data[4024]=8'b01100010;
   assign rom_data[4025]=8'b10000010;
   assign rom_data[4026]=8'b01100010;
   assign rom_data[4027]=8'b10000011;
   assign rom_data[4028]=8'b01100010;
   assign rom_data[4029]=8'b10000100;
   assign rom_data[4030]=8'b01100010;
   assign rom_data[4031]=8'b10000101;
   assign rom_data[4032]=8'b01100010;
   assign rom_data[4033]=8'b10000110;
   assign rom_data[4034]=8'b01100010;
   assign rom_data[4035]=8'b10000110;
   assign rom_data[4036]=8'b01100010;
   assign rom_data[4037]=8'b10000111;
   assign rom_data[4038]=8'b01100010;
   assign rom_data[4039]=8'b10001000;
   assign rom_data[4040]=8'b01100010;
   assign rom_data[4041]=8'b10001000;
   assign rom_data[4042]=8'b01100010;
   assign rom_data[4043]=8'b10001001;
   assign rom_data[4044]=8'b01100010;
   assign rom_data[4045]=8'b10001001;
   assign rom_data[4046]=8'b01100010;
   assign rom_data[4047]=8'b10001001;
   assign rom_data[4048]=8'b01100010;
   assign rom_data[4049]=8'b10001010;
   assign rom_data[4050]=8'b01100010;
   assign rom_data[4051]=8'b10001010;
   assign rom_data[4052]=8'b01100010;
   assign rom_data[4053]=8'b10001010;
   assign rom_data[4054]=8'b01100010;
   assign rom_data[4055]=8'b10001010;
   assign rom_data[4056]=8'b01100010;
   assign rom_data[4057]=8'b10001010;
   assign rom_data[4058]=8'b01100010;
   assign rom_data[4059]=8'b10001001;
   assign rom_data[4060]=8'b01100010;
   assign rom_data[4061]=8'b10001001;
   assign rom_data[4062]=8'b01100010;
   assign rom_data[4063]=8'b10001001;
   assign rom_data[4064]=8'b01100010;
   assign rom_data[4065]=8'b10001000;
   assign rom_data[4066]=8'b01100010;
   assign rom_data[4067]=8'b10001000;
   assign rom_data[4068]=8'b01100010;
   assign rom_data[4069]=8'b10000111;
   assign rom_data[4070]=8'b01100010;
   assign rom_data[4071]=8'b10000111;
   assign rom_data[4072]=8'b01100010;
   assign rom_data[4073]=8'b10000110;
   assign rom_data[4074]=8'b01100010;
   assign rom_data[4075]=8'b10000101;
   assign rom_data[4076]=8'b01100011;
   assign rom_data[4077]=8'b10000100;
   assign rom_data[4078]=8'b01100011;
   assign rom_data[4079]=8'b10000011;
   assign rom_data[4080]=8'b01100011;
   assign rom_data[4081]=8'b10000011;
   assign rom_data[4082]=8'b01100011;
   assign rom_data[4083]=8'b10000010;
   assign rom_data[4084]=8'b01100011;
   assign rom_data[4085]=8'b10000001;
   assign rom_data[4086]=8'b01100011;
   assign rom_data[4087]=8'b10000000;
   assign rom_data[4088]=8'b01100011;
   assign rom_data[4089]=8'b01111110;
   assign rom_data[4090]=8'b01100011;
   assign rom_data[4091]=8'b01111101;
   assign rom_data[4092]=8'b01100011;
   assign rom_data[4093]=8'b01111100;
   assign rom_data[4094]=8'b01100011;
   assign rom_data[4095]=8'b01111011;
   assign rom_data[4096]=8'b01100011;
   assign rom_data[4097]=8'b01111010;
   assign rom_data[4098]=8'b01100011;
   assign rom_data[4099]=8'b01111001;
   assign rom_data[4100]=8'b01100011;
   assign rom_data[4101]=8'b01110111;
   assign rom_data[4102]=8'b01100011;
   assign rom_data[4103]=8'b01110110;
   assign rom_data[4104]=8'b01100011;
   assign rom_data[4105]=8'b01110101;
   assign rom_data[4106]=8'b01100011;
   assign rom_data[4107]=8'b01110100;
   assign rom_data[4108]=8'b01100011;
   assign rom_data[4109]=8'b01110010;
   assign rom_data[4110]=8'b01100011;
   assign rom_data[4111]=8'b01110001;
   assign rom_data[4112]=8'b01100011;
   assign rom_data[4113]=8'b01110000;
   assign rom_data[4114]=8'b01100011;
   assign rom_data[4115]=8'b01101110;
   assign rom_data[4116]=8'b01100011;
   assign rom_data[4117]=8'b01101101;
   assign rom_data[4118]=8'b01100011;
   assign rom_data[4119]=8'b01101100;
   assign rom_data[4120]=8'b01100011;
   assign rom_data[4121]=8'b01101010;
   assign rom_data[4122]=8'b01100011;
   assign rom_data[4123]=8'b01101001;
   assign rom_data[4124]=8'b01100011;
   assign rom_data[4125]=8'b01100111;
   assign rom_data[4126]=8'b01100011;
   assign rom_data[4127]=8'b01100110;
   assign rom_data[4128]=8'b01100011;
   assign rom_data[4129]=8'b01100101;
   assign rom_data[4130]=8'b01100011;
   assign rom_data[4131]=8'b01100011;
   assign rom_data[4132]=8'b01100011;
   assign rom_data[4133]=8'b01100010;
   assign rom_data[4134]=8'b01100011;
   assign rom_data[4135]=8'b01100001;
   assign rom_data[4136]=8'b01100011;
   assign rom_data[4137]=8'b01011111;
   assign rom_data[4138]=8'b01100011;
   assign rom_data[4139]=8'b01011110;
   assign rom_data[4140]=8'b01100011;
   assign rom_data[4141]=8'b01011100;
   assign rom_data[4142]=8'b01100011;
   assign rom_data[4143]=8'b01011011;
   assign rom_data[4144]=8'b01100011;
   assign rom_data[4145]=8'b01011001;
   assign rom_data[4146]=8'b01100011;
   assign rom_data[4147]=8'b01011000;
   assign rom_data[4148]=8'b01100011;
   assign rom_data[4149]=8'b01010111;
   assign rom_data[4150]=8'b01100011;
   assign rom_data[4151]=8'b01010101;
   assign rom_data[4152]=8'b01100011;
   assign rom_data[4153]=8'b01010100;
   assign rom_data[4154]=8'b01100011;
   assign rom_data[4155]=8'b01010010;
   assign rom_data[4156]=8'b01100011;
   assign rom_data[4157]=8'b01010001;
   assign rom_data[4158]=8'b01100100;
   assign rom_data[4159]=8'b01010000;
   assign rom_data[4160]=8'b01100100;
   assign rom_data[4161]=8'b01001110;
   assign rom_data[4162]=8'b01100100;
   assign rom_data[4163]=8'b01001101;
   assign rom_data[4164]=8'b01100100;
   assign rom_data[4165]=8'b01001100;
   assign rom_data[4166]=8'b01100100;
   assign rom_data[4167]=8'b01001010;
   assign rom_data[4168]=8'b01100100;
   assign rom_data[4169]=8'b01001001;
   assign rom_data[4170]=8'b01100100;
   assign rom_data[4171]=8'b01001000;
   assign rom_data[4172]=8'b01100100;
   assign rom_data[4173]=8'b01000110;
   assign rom_data[4174]=8'b01100100;
   assign rom_data[4175]=8'b01000101;
   assign rom_data[4176]=8'b01100100;
   assign rom_data[4177]=8'b01000100;
   assign rom_data[4178]=8'b01100100;
   assign rom_data[4179]=8'b01000010;
   assign rom_data[4180]=8'b01100100;
   assign rom_data[4181]=8'b01000001;
   assign rom_data[4182]=8'b01100100;
   assign rom_data[4183]=8'b01000000;
   assign rom_data[4184]=8'b01100100;
   assign rom_data[4185]=8'b00111111;
   assign rom_data[4186]=8'b01100100;
   assign rom_data[4187]=8'b00111101;
   assign rom_data[4188]=8'b01100100;
   assign rom_data[4189]=8'b00111100;
   assign rom_data[4190]=8'b01100100;
   assign rom_data[4191]=8'b00111011;
   assign rom_data[4192]=8'b01100100;
   assign rom_data[4193]=8'b00111010;
   assign rom_data[4194]=8'b01100100;
   assign rom_data[4195]=8'b00111001;
   assign rom_data[4196]=8'b01100100;
   assign rom_data[4197]=8'b00111000;
   assign rom_data[4198]=8'b01100100;
   assign rom_data[4199]=8'b00110110;
   assign rom_data[4200]=8'b01100100;
   assign rom_data[4201]=8'b00110101;
   assign rom_data[4202]=8'b01100100;
   assign rom_data[4203]=8'b00110100;
   assign rom_data[4204]=8'b01100100;
   assign rom_data[4205]=8'b00110011;
   assign rom_data[4206]=8'b01100100;
   assign rom_data[4207]=8'b00110011;
   assign rom_data[4208]=8'b01100100;
   assign rom_data[4209]=8'b00110010;
   assign rom_data[4210]=8'b01100100;
   assign rom_data[4211]=8'b00110001;
   assign rom_data[4212]=8'b01100100;
   assign rom_data[4213]=8'b00110000;
   assign rom_data[4214]=8'b01100100;
   assign rom_data[4215]=8'b00101111;
   assign rom_data[4216]=8'b01100100;
   assign rom_data[4217]=8'b00101111;
   assign rom_data[4218]=8'b01100100;
   assign rom_data[4219]=8'b00101110;
   assign rom_data[4220]=8'b01100100;
   assign rom_data[4221]=8'b00101110;
   assign rom_data[4222]=8'b01100100;
   assign rom_data[4223]=8'b00101101;
   assign rom_data[4224]=8'b01100100;
   assign rom_data[4225]=8'b00101101;
   assign rom_data[4226]=8'b01100100;
   assign rom_data[4227]=8'b00101100;
   assign rom_data[4228]=8'b01100100;
   assign rom_data[4229]=8'b00101100;
   assign rom_data[4230]=8'b01100100;
   assign rom_data[4231]=8'b00101100;
   assign rom_data[4232]=8'b01100101;
   assign rom_data[4233]=8'b00101100;
   assign rom_data[4234]=8'b01100101;
   assign rom_data[4235]=8'b00101100;
   assign rom_data[4236]=8'b01100101;
   assign rom_data[4237]=8'b00101100;
   assign rom_data[4238]=8'b01100101;
   assign rom_data[4239]=8'b00101100;
   assign rom_data[4240]=8'b01100101;
   assign rom_data[4241]=8'b00101101;
   assign rom_data[4242]=8'b01100101;
   assign rom_data[4243]=8'b00101101;
   assign rom_data[4244]=8'b01100101;
   assign rom_data[4245]=8'b00101101;
   assign rom_data[4246]=8'b01100101;
   assign rom_data[4247]=8'b00101110;
   assign rom_data[4248]=8'b01100101;
   assign rom_data[4249]=8'b00101111;
   assign rom_data[4250]=8'b01100101;
   assign rom_data[4251]=8'b00101111;
   assign rom_data[4252]=8'b01100101;
   assign rom_data[4253]=8'b00110000;
   assign rom_data[4254]=8'b01100101;
   assign rom_data[4255]=8'b00110001;
   assign rom_data[4256]=8'b01100101;
   assign rom_data[4257]=8'b00110001;
   assign rom_data[4258]=8'b01100101;
   assign rom_data[4259]=8'b00110010;
   assign rom_data[4260]=8'b01100101;
   assign rom_data[4261]=8'b00110011;
   assign rom_data[4262]=8'b01100101;
   assign rom_data[4263]=8'b00110100;
   assign rom_data[4264]=8'b01100101;
   assign rom_data[4265]=8'b00110101;
   assign rom_data[4266]=8'b01100101;
   assign rom_data[4267]=8'b00110110;
   assign rom_data[4268]=8'b01100101;
   assign rom_data[4269]=8'b00110111;
   assign rom_data[4270]=8'b01100101;
   assign rom_data[4271]=8'b00111000;
   assign rom_data[4272]=8'b01100101;
   assign rom_data[4273]=8'b00111010;
   assign rom_data[4274]=8'b01100101;
   assign rom_data[4275]=8'b00111011;
   assign rom_data[4276]=8'b01100101;
   assign rom_data[4277]=8'b00111100;
   assign rom_data[4278]=8'b01100101;
   assign rom_data[4279]=8'b00111101;
   assign rom_data[4280]=8'b01100101;
   assign rom_data[4281]=8'b00111110;
   assign rom_data[4282]=8'b01100101;
   assign rom_data[4283]=8'b01000000;
   assign rom_data[4284]=8'b01100101;
   assign rom_data[4285]=8'b01000001;
   assign rom_data[4286]=8'b01100101;
   assign rom_data[4287]=8'b01000010;
   assign rom_data[4288]=8'b01100101;
   assign rom_data[4289]=8'b01000100;
   assign rom_data[4290]=8'b01100101;
   assign rom_data[4291]=8'b01000101;
   assign rom_data[4292]=8'b01100101;
   assign rom_data[4293]=8'b01000110;
   assign rom_data[4294]=8'b01100101;
   assign rom_data[4295]=8'b01001000;
   assign rom_data[4296]=8'b01100101;
   assign rom_data[4297]=8'b01001001;
   assign rom_data[4298]=8'b01100101;
   assign rom_data[4299]=8'b01001010;
   assign rom_data[4300]=8'b01100101;
   assign rom_data[4301]=8'b01001100;
   assign rom_data[4302]=8'b01100110;
   assign rom_data[4303]=8'b01001101;
   assign rom_data[4304]=8'b01100110;
   assign rom_data[4305]=8'b01001110;
   assign rom_data[4306]=8'b01100110;
   assign rom_data[4307]=8'b01010000;
   assign rom_data[4308]=8'b01100110;
   assign rom_data[4309]=8'b01010001;
   assign rom_data[4310]=8'b01100110;
   assign rom_data[4311]=8'b01010011;
   assign rom_data[4312]=8'b01100110;
   assign rom_data[4313]=8'b01010100;
   assign rom_data[4314]=8'b01100110;
   assign rom_data[4315]=8'b01010101;
   assign rom_data[4316]=8'b01100110;
   assign rom_data[4317]=8'b01010111;
   assign rom_data[4318]=8'b01100110;
   assign rom_data[4319]=8'b01011000;
   assign rom_data[4320]=8'b01100110;
   assign rom_data[4321]=8'b01011010;
   assign rom_data[4322]=8'b01100110;
   assign rom_data[4323]=8'b01011011;
   assign rom_data[4324]=8'b01100110;
   assign rom_data[4325]=8'b01011100;
   assign rom_data[4326]=8'b01100110;
   assign rom_data[4327]=8'b01011110;
   assign rom_data[4328]=8'b01100110;
   assign rom_data[4329]=8'b01011111;
   assign rom_data[4330]=8'b01100110;
   assign rom_data[4331]=8'b01100001;
   assign rom_data[4332]=8'b01100110;
   assign rom_data[4333]=8'b01100010;
   assign rom_data[4334]=8'b01100110;
   assign rom_data[4335]=8'b01100011;
   assign rom_data[4336]=8'b01100110;
   assign rom_data[4337]=8'b01100101;
   assign rom_data[4338]=8'b01100110;
   assign rom_data[4339]=8'b01100110;
   assign rom_data[4340]=8'b01100110;
   assign rom_data[4341]=8'b01101000;
   assign rom_data[4342]=8'b01100110;
   assign rom_data[4343]=8'b01101001;
   assign rom_data[4344]=8'b01100110;
   assign rom_data[4345]=8'b01101010;
   assign rom_data[4346]=8'b01100110;
   assign rom_data[4347]=8'b01101100;
   assign rom_data[4348]=8'b01100110;
   assign rom_data[4349]=8'b01101101;
   assign rom_data[4350]=8'b01100110;
   assign rom_data[4351]=8'b01101110;
   assign rom_data[4352]=8'b01100110;
   assign rom_data[4353]=8'b01110000;
   assign rom_data[4354]=8'b01100110;
   assign rom_data[4355]=8'b01110001;
   assign rom_data[4356]=8'b01100110;
   assign rom_data[4357]=8'b01110010;
   assign rom_data[4358]=8'b01100110;
   assign rom_data[4359]=8'b01110100;
   assign rom_data[4360]=8'b01100110;
   assign rom_data[4361]=8'b01110101;
   assign rom_data[4362]=8'b01100110;
   assign rom_data[4363]=8'b01110110;
   assign rom_data[4364]=8'b01100110;
   assign rom_data[4365]=8'b01110111;
   assign rom_data[4366]=8'b01100110;
   assign rom_data[4367]=8'b01111001;
   assign rom_data[4368]=8'b01100110;
   assign rom_data[4369]=8'b01111010;
   assign rom_data[4370]=8'b01100110;
   assign rom_data[4371]=8'b01111011;
   assign rom_data[4372]=8'b01100110;
   assign rom_data[4373]=8'b01111100;
   assign rom_data[4374]=8'b01100110;
   assign rom_data[4375]=8'b01111101;
   assign rom_data[4376]=8'b01100110;
   assign rom_data[4377]=8'b01111110;
   assign rom_data[4378]=8'b01100110;
   assign rom_data[4379]=8'b01111111;
   assign rom_data[4380]=8'b01100110;
   assign rom_data[4381]=8'b10000000;
   assign rom_data[4382]=8'b01100110;
   assign rom_data[4383]=8'b10000001;
   assign rom_data[4384]=8'b01100111;
   assign rom_data[4385]=8'b10000010;
   assign rom_data[4386]=8'b01100111;
   assign rom_data[4387]=8'b10000011;
   assign rom_data[4388]=8'b01100111;
   assign rom_data[4389]=8'b10000100;
   assign rom_data[4390]=8'b01100111;
   assign rom_data[4391]=8'b10000101;
   assign rom_data[4392]=8'b01100111;
   assign rom_data[4393]=8'b10000110;
   assign rom_data[4394]=8'b01100111;
   assign rom_data[4395]=8'b10000110;
   assign rom_data[4396]=8'b01100111;
   assign rom_data[4397]=8'b10000111;
   assign rom_data[4398]=8'b01100111;
   assign rom_data[4399]=8'b10001000;
   assign rom_data[4400]=8'b01100111;
   assign rom_data[4401]=8'b10001000;
   assign rom_data[4402]=8'b01100111;
   assign rom_data[4403]=8'b10001001;
   assign rom_data[4404]=8'b01100111;
   assign rom_data[4405]=8'b10001001;
   assign rom_data[4406]=8'b01100111;
   assign rom_data[4407]=8'b10001001;
   assign rom_data[4408]=8'b01100111;
   assign rom_data[4409]=8'b10001010;
   assign rom_data[4410]=8'b01100111;
   assign rom_data[4411]=8'b10001010;
   assign rom_data[4412]=8'b01100111;
   assign rom_data[4413]=8'b10001010;
   assign rom_data[4414]=8'b01100111;
   assign rom_data[4415]=8'b10001010;
   assign rom_data[4416]=8'b01100111;
   assign rom_data[4417]=8'b10001010;
   assign rom_data[4418]=8'b01100111;
   assign rom_data[4419]=8'b10001001;
   assign rom_data[4420]=8'b01100111;
   assign rom_data[4421]=8'b10001001;
   assign rom_data[4422]=8'b01100111;
   assign rom_data[4423]=8'b10001001;
   assign rom_data[4424]=8'b01100111;
   assign rom_data[4425]=8'b10001000;
   assign rom_data[4426]=8'b01100111;
   assign rom_data[4427]=8'b10001000;
   assign rom_data[4428]=8'b01100111;
   assign rom_data[4429]=8'b10000111;
   assign rom_data[4430]=8'b01100111;
   assign rom_data[4431]=8'b10000111;
   assign rom_data[4432]=8'b01100111;
   assign rom_data[4433]=8'b10000110;
   assign rom_data[4434]=8'b01100111;
   assign rom_data[4435]=8'b10000101;
   assign rom_data[4436]=8'b01100111;
   assign rom_data[4437]=8'b10000100;
   assign rom_data[4438]=8'b01100111;
   assign rom_data[4439]=8'b10000011;
   assign rom_data[4440]=8'b01100111;
   assign rom_data[4441]=8'b10000011;
   assign rom_data[4442]=8'b01100111;
   assign rom_data[4443]=8'b10000010;
   assign rom_data[4444]=8'b01100111;
   assign rom_data[4445]=8'b10000001;
   assign rom_data[4446]=8'b01100111;
   assign rom_data[4447]=8'b10000000;
   assign rom_data[4448]=8'b01100111;
   assign rom_data[4449]=8'b01111110;
   assign rom_data[4450]=8'b01101000;
   assign rom_data[4451]=8'b01111101;
   assign rom_data[4452]=8'b01101000;
   assign rom_data[4453]=8'b01111100;
   assign rom_data[4454]=8'b01101000;
   assign rom_data[4455]=8'b01111011;
   assign rom_data[4456]=8'b01101000;
   assign rom_data[4457]=8'b01111010;
   assign rom_data[4458]=8'b01101000;
   assign rom_data[4459]=8'b01111001;
   assign rom_data[4460]=8'b01101000;
   assign rom_data[4461]=8'b01110111;
   assign rom_data[4462]=8'b01101000;
   assign rom_data[4463]=8'b01110110;
   assign rom_data[4464]=8'b01101000;
   assign rom_data[4465]=8'b01110101;
   assign rom_data[4466]=8'b01101000;
   assign rom_data[4467]=8'b01110100;
   assign rom_data[4468]=8'b01101000;
   assign rom_data[4469]=8'b01110010;
   assign rom_data[4470]=8'b01101000;
   assign rom_data[4471]=8'b01110001;
   assign rom_data[4472]=8'b01101000;
   assign rom_data[4473]=8'b01110000;
   assign rom_data[4474]=8'b01101000;
   assign rom_data[4475]=8'b01101110;
   assign rom_data[4476]=8'b01101000;
   assign rom_data[4477]=8'b01101101;
   assign rom_data[4478]=8'b01101000;
   assign rom_data[4479]=8'b01101100;
   assign rom_data[4480]=8'b01101000;
   assign rom_data[4481]=8'b01101010;
   assign rom_data[4482]=8'b01101000;
   assign rom_data[4483]=8'b01101001;
   assign rom_data[4484]=8'b01101000;
   assign rom_data[4485]=8'b01100111;
   assign rom_data[4486]=8'b01101000;
   assign rom_data[4487]=8'b01100110;
   assign rom_data[4488]=8'b01101000;
   assign rom_data[4489]=8'b01100101;
   assign rom_data[4490]=8'b01101000;
   assign rom_data[4491]=8'b01100011;
   assign rom_data[4492]=8'b01101000;
   assign rom_data[4493]=8'b01100010;
   assign rom_data[4494]=8'b01101000;
   assign rom_data[4495]=8'b01100001;
   assign rom_data[4496]=8'b01101000;
   assign rom_data[4497]=8'b01011111;
   assign rom_data[4498]=8'b01101000;
   assign rom_data[4499]=8'b01011110;
   assign rom_data[4500]=8'b01101000;
   assign rom_data[4501]=8'b01011100;
   assign rom_data[4502]=8'b01101000;
   assign rom_data[4503]=8'b01011011;
   assign rom_data[4504]=8'b01101000;
   assign rom_data[4505]=8'b01011001;
   assign rom_data[4506]=8'b01101000;
   assign rom_data[4507]=8'b01011000;
   assign rom_data[4508]=8'b01101000;
   assign rom_data[4509]=8'b01010111;
   assign rom_data[4510]=8'b01101000;
   assign rom_data[4511]=8'b01010101;
   assign rom_data[4512]=8'b01101000;
   assign rom_data[4513]=8'b01010100;
   assign rom_data[4514]=8'b01101000;
   assign rom_data[4515]=8'b01010010;
   assign rom_data[4516]=8'b01101000;
   assign rom_data[4517]=8'b01010001;
   assign rom_data[4518]=8'b01101000;
   assign rom_data[4519]=8'b01010000;
   assign rom_data[4520]=8'b01101000;
   assign rom_data[4521]=8'b01001110;
   assign rom_data[4522]=8'b01101000;
   assign rom_data[4523]=8'b01001101;
   assign rom_data[4524]=8'b01101000;
   assign rom_data[4525]=8'b01001100;
   assign rom_data[4526]=8'b01101000;
   assign rom_data[4527]=8'b01001010;
   assign rom_data[4528]=8'b01101000;
   assign rom_data[4529]=8'b01001001;
   assign rom_data[4530]=8'b01101000;
   assign rom_data[4531]=8'b01001000;
   assign rom_data[4532]=8'b01101000;
   assign rom_data[4533]=8'b01000110;
   assign rom_data[4534]=8'b01101001;
   assign rom_data[4535]=8'b01000101;
   assign rom_data[4536]=8'b01101001;
   assign rom_data[4537]=8'b01000100;
   assign rom_data[4538]=8'b01101001;
   assign rom_data[4539]=8'b01000010;
   assign rom_data[4540]=8'b01101001;
   assign rom_data[4541]=8'b01000001;
   assign rom_data[4542]=8'b01101001;
   assign rom_data[4543]=8'b01000000;
   assign rom_data[4544]=8'b01101001;
   assign rom_data[4545]=8'b00111111;
   assign rom_data[4546]=8'b01101001;
   assign rom_data[4547]=8'b00111101;
   assign rom_data[4548]=8'b01101001;
   assign rom_data[4549]=8'b00111100;
   assign rom_data[4550]=8'b01101001;
   assign rom_data[4551]=8'b00111011;
   assign rom_data[4552]=8'b01101001;
   assign rom_data[4553]=8'b00111010;
   assign rom_data[4554]=8'b01101001;
   assign rom_data[4555]=8'b00111001;
   assign rom_data[4556]=8'b01101001;
   assign rom_data[4557]=8'b00111000;
   assign rom_data[4558]=8'b01101001;
   assign rom_data[4559]=8'b00110110;
   assign rom_data[4560]=8'b01101001;
   assign rom_data[4561]=8'b00110101;
   assign rom_data[4562]=8'b01101001;
   assign rom_data[4563]=8'b00110100;
   assign rom_data[4564]=8'b01101001;
   assign rom_data[4565]=8'b00110011;
   assign rom_data[4566]=8'b01101001;
   assign rom_data[4567]=8'b00110011;
   assign rom_data[4568]=8'b01101001;
   assign rom_data[4569]=8'b00110010;
   assign rom_data[4570]=8'b01101001;
   assign rom_data[4571]=8'b00110001;
   assign rom_data[4572]=8'b01101001;
   assign rom_data[4573]=8'b00110000;
   assign rom_data[4574]=8'b01101001;
   assign rom_data[4575]=8'b00101111;
   assign rom_data[4576]=8'b01101001;
   assign rom_data[4577]=8'b00101111;
   assign rom_data[4578]=8'b01101001;
   assign rom_data[4579]=8'b00101110;
   assign rom_data[4580]=8'b01101001;
   assign rom_data[4581]=8'b00101110;
   assign rom_data[4582]=8'b01101001;
   assign rom_data[4583]=8'b00101101;
   assign rom_data[4584]=8'b01101001;
   assign rom_data[4585]=8'b00101101;
   assign rom_data[4586]=8'b01101001;
   assign rom_data[4587]=8'b00101100;
   assign rom_data[4588]=8'b01101001;
   assign rom_data[4589]=8'b00101100;
   assign rom_data[4590]=8'b01101001;
   assign rom_data[4591]=8'b00101100;
   assign rom_data[4592]=8'b01101001;
   assign rom_data[4593]=8'b00101100;
   assign rom_data[4594]=8'b01101001;
   assign rom_data[4595]=8'b00101100;
   assign rom_data[4596]=8'b01101001;
   assign rom_data[4597]=8'b00101100;
   assign rom_data[4598]=8'b01101001;
   assign rom_data[4599]=8'b00101100;
   assign rom_data[4600]=8'b01101001;
   assign rom_data[4601]=8'b00101101;
   assign rom_data[4602]=8'b01101010;
   assign rom_data[4603]=8'b00101101;
   assign rom_data[4604]=8'b01101010;
   assign rom_data[4605]=8'b00101101;
   assign rom_data[4606]=8'b01101010;
   assign rom_data[4607]=8'b00101110;
   assign rom_data[4608]=8'b01101010;
   assign rom_data[4609]=8'b00101111;
   assign rom_data[4610]=8'b01101010;
   assign rom_data[4611]=8'b00101111;
   assign rom_data[4612]=8'b01101010;
   assign rom_data[4613]=8'b00110000;
   assign rom_data[4614]=8'b01101010;
   assign rom_data[4615]=8'b00110001;
   assign rom_data[4616]=8'b01101010;
   assign rom_data[4617]=8'b00110001;
   assign rom_data[4618]=8'b01101010;
   assign rom_data[4619]=8'b00110010;
   assign rom_data[4620]=8'b01101010;
   assign rom_data[4621]=8'b00110011;
   assign rom_data[4622]=8'b01101010;
   assign rom_data[4623]=8'b00110100;
   assign rom_data[4624]=8'b01101010;
   assign rom_data[4625]=8'b00110101;
   assign rom_data[4626]=8'b01101010;
   assign rom_data[4627]=8'b00110110;
   assign rom_data[4628]=8'b01101010;
   assign rom_data[4629]=8'b00110111;
   assign rom_data[4630]=8'b01101010;
   assign rom_data[4631]=8'b00111000;
   assign rom_data[4632]=8'b01101010;
   assign rom_data[4633]=8'b00111010;
   assign rom_data[4634]=8'b01101010;
   assign rom_data[4635]=8'b00111011;
   assign rom_data[4636]=8'b01101010;
   assign rom_data[4637]=8'b00111100;
   assign rom_data[4638]=8'b01101010;
   assign rom_data[4639]=8'b00111101;
   assign rom_data[4640]=8'b01101010;
   assign rom_data[4641]=8'b00111110;
   assign rom_data[4642]=8'b01101010;
   assign rom_data[4643]=8'b01000000;
   assign rom_data[4644]=8'b01101010;
   assign rom_data[4645]=8'b01000001;
   assign rom_data[4646]=8'b01101010;
   assign rom_data[4647]=8'b01000010;
   assign rom_data[4648]=8'b01101010;
   assign rom_data[4649]=8'b01000100;
   assign rom_data[4650]=8'b01101010;
   assign rom_data[4651]=8'b01000101;
   assign rom_data[4652]=8'b01101010;
   assign rom_data[4653]=8'b01000110;
   assign rom_data[4654]=8'b01101010;
   assign rom_data[4655]=8'b01001000;
   assign rom_data[4656]=8'b01101010;
   assign rom_data[4657]=8'b01001001;
   assign rom_data[4658]=8'b01101010;
   assign rom_data[4659]=8'b01001010;
   assign rom_data[4660]=8'b01101010;
   assign rom_data[4661]=8'b01001100;
   assign rom_data[4662]=8'b01101010;
   assign rom_data[4663]=8'b01001101;
   assign rom_data[4664]=8'b01101010;
   assign rom_data[4665]=8'b01001110;
   assign rom_data[4666]=8'b01101010;
   assign rom_data[4667]=8'b01010000;
   assign rom_data[4668]=8'b01101010;
   assign rom_data[4669]=8'b01010001;
   assign rom_data[4670]=8'b01101010;
   assign rom_data[4671]=8'b01010011;
   assign rom_data[4672]=8'b01101010;
   assign rom_data[4673]=8'b01010100;
   assign rom_data[4674]=8'b01101010;
   assign rom_data[4675]=8'b01010101;
   assign rom_data[4676]=8'b01101010;
   assign rom_data[4677]=8'b01010111;
   assign rom_data[4678]=8'b01101011;
   assign rom_data[4679]=8'b01011000;
   assign rom_data[4680]=8'b01101011;
   assign rom_data[4681]=8'b01011010;
   assign rom_data[4682]=8'b01101011;
   assign rom_data[4683]=8'b01011011;
   assign rom_data[4684]=8'b01101011;
   assign rom_data[4685]=8'b01011100;
   assign rom_data[4686]=8'b01101011;
   assign rom_data[4687]=8'b01011110;
   assign rom_data[4688]=8'b01101011;
   assign rom_data[4689]=8'b01011111;
   assign rom_data[4690]=8'b01101011;
   assign rom_data[4691]=8'b01100001;
   assign rom_data[4692]=8'b01101011;
   assign rom_data[4693]=8'b01100010;
   assign rom_data[4694]=8'b01101011;
   assign rom_data[4695]=8'b01100011;
   assign rom_data[4696]=8'b01101011;
   assign rom_data[4697]=8'b01100101;
   assign rom_data[4698]=8'b01101011;
   assign rom_data[4699]=8'b01100110;
   assign rom_data[4700]=8'b01101011;
   assign rom_data[4701]=8'b01101000;
   assign rom_data[4702]=8'b01101011;
   assign rom_data[4703]=8'b01101001;
   assign rom_data[4704]=8'b01101011;
   assign rom_data[4705]=8'b01101010;
   assign rom_data[4706]=8'b01101011;
   assign rom_data[4707]=8'b01101100;
   assign rom_data[4708]=8'b01101011;
   assign rom_data[4709]=8'b01101101;
   assign rom_data[4710]=8'b01101011;
   assign rom_data[4711]=8'b01101110;
   assign rom_data[4712]=8'b01101011;
   assign rom_data[4713]=8'b01110000;
   assign rom_data[4714]=8'b01101011;
   assign rom_data[4715]=8'b01110001;
   assign rom_data[4716]=8'b01101011;
   assign rom_data[4717]=8'b01110010;
   assign rom_data[4718]=8'b01101011;
   assign rom_data[4719]=8'b01110100;
   assign rom_data[4720]=8'b01101011;
   assign rom_data[4721]=8'b01110101;
   assign rom_data[4722]=8'b01101011;
   assign rom_data[4723]=8'b01110110;
   assign rom_data[4724]=8'b01101011;
   assign rom_data[4725]=8'b01110111;
   assign rom_data[4726]=8'b01101011;
   assign rom_data[4727]=8'b01111001;
   assign rom_data[4728]=8'b01101011;
   assign rom_data[4729]=8'b01111010;
   assign rom_data[4730]=8'b01101011;
   assign rom_data[4731]=8'b01111011;
   assign rom_data[4732]=8'b01101011;
   assign rom_data[4733]=8'b01111100;
   assign rom_data[4734]=8'b01101011;
   assign rom_data[4735]=8'b01111101;
   assign rom_data[4736]=8'b01101011;
   assign rom_data[4737]=8'b01111110;
   assign rom_data[4738]=8'b01101011;
   assign rom_data[4739]=8'b01111111;
   assign rom_data[4740]=8'b01101011;
   assign rom_data[4741]=8'b10000000;
   assign rom_data[4742]=8'b01101011;
   assign rom_data[4743]=8'b10000001;
   assign rom_data[4744]=8'b01101011;
   assign rom_data[4745]=8'b10000010;
   assign rom_data[4746]=8'b01101011;
   assign rom_data[4747]=8'b10000011;
   assign rom_data[4748]=8'b01101011;
   assign rom_data[4749]=8'b10000100;
   assign rom_data[4750]=8'b01101011;
   assign rom_data[4751]=8'b10000101;
   assign rom_data[4752]=8'b01101011;
   assign rom_data[4753]=8'b10000110;
   assign rom_data[4754]=8'b01101011;
   assign rom_data[4755]=8'b10000110;
   assign rom_data[4756]=8'b01101011;
   assign rom_data[4757]=8'b10000111;
   assign rom_data[4758]=8'b01101100;
   assign rom_data[4759]=8'b10001000;
   assign rom_data[4760]=8'b01101100;
   assign rom_data[4761]=8'b10001000;
   assign rom_data[4762]=8'b01101100;
   assign rom_data[4763]=8'b10001001;
   assign rom_data[4764]=8'b01101100;
   assign rom_data[4765]=8'b10001001;
   assign rom_data[4766]=8'b01101100;
   assign rom_data[4767]=8'b10001001;
   assign rom_data[4768]=8'b01101100;
   assign rom_data[4769]=8'b10001010;
   assign rom_data[4770]=8'b01101100;
   assign rom_data[4771]=8'b10001010;
   assign rom_data[4772]=8'b01101100;
   assign rom_data[4773]=8'b10001010;
   assign rom_data[4774]=8'b01101100;
   assign rom_data[4775]=8'b10001010;
   assign rom_data[4776]=8'b01101100;
   assign rom_data[4777]=8'b10001010;
   assign rom_data[4778]=8'b01101100;
   assign rom_data[4779]=8'b10001001;
   assign rom_data[4780]=8'b01101100;
   assign rom_data[4781]=8'b10001001;
   assign rom_data[4782]=8'b01101100;
   assign rom_data[4783]=8'b10001001;
   assign rom_data[4784]=8'b01101100;
   assign rom_data[4785]=8'b10001000;
   assign rom_data[4786]=8'b01101100;
   assign rom_data[4787]=8'b10001000;
   assign rom_data[4788]=8'b01101100;
   assign rom_data[4789]=8'b10000111;
   assign rom_data[4790]=8'b01101100;
   assign rom_data[4791]=8'b10000111;
   assign rom_data[4792]=8'b01101100;
   assign rom_data[4793]=8'b10000110;
   assign rom_data[4794]=8'b01101100;
   assign rom_data[4795]=8'b10000101;
   assign rom_data[4796]=8'b01101100;
   assign rom_data[4797]=8'b10000100;
   assign rom_data[4798]=8'b01101100;
   assign rom_data[4799]=8'b10000011;
   assign rom_data[4800]=8'b01101100;
   assign rom_data[4801]=8'b10000011;
   assign rom_data[4802]=8'b01101100;
   assign rom_data[4803]=8'b10000010;
   assign rom_data[4804]=8'b01101100;
   assign rom_data[4805]=8'b10000001;
   assign rom_data[4806]=8'b01101100;
   assign rom_data[4807]=8'b10000000;
   assign rom_data[4808]=8'b01101100;
   assign rom_data[4809]=8'b01111110;
   assign rom_data[4810]=8'b01101100;
   assign rom_data[4811]=8'b01111101;
   assign rom_data[4812]=8'b01101100;
   assign rom_data[4813]=8'b01111100;
   assign rom_data[4814]=8'b01101100;
   assign rom_data[4815]=8'b01111011;
   assign rom_data[4816]=8'b01101100;
   assign rom_data[4817]=8'b01111010;
   assign rom_data[4818]=8'b01101100;
   assign rom_data[4819]=8'b01111001;
   assign rom_data[4820]=8'b01101100;
   assign rom_data[4821]=8'b01110111;
   assign rom_data[4822]=8'b01101100;
   assign rom_data[4823]=8'b01110110;
   assign rom_data[4824]=8'b01101101;
   assign rom_data[4825]=8'b01110101;
   assign rom_data[4826]=8'b01101101;
   assign rom_data[4827]=8'b01110100;
   assign rom_data[4828]=8'b01101101;
   assign rom_data[4829]=8'b01110010;
   assign rom_data[4830]=8'b01101101;
   assign rom_data[4831]=8'b01110001;
   assign rom_data[4832]=8'b01101101;
   assign rom_data[4833]=8'b01110000;
   assign rom_data[4834]=8'b01101101;
   assign rom_data[4835]=8'b01101110;
   assign rom_data[4836]=8'b01101101;
   assign rom_data[4837]=8'b01101101;
   assign rom_data[4838]=8'b01101101;
   assign rom_data[4839]=8'b01101100;
   assign rom_data[4840]=8'b01101101;
   assign rom_data[4841]=8'b01101010;
   assign rom_data[4842]=8'b01101101;
   assign rom_data[4843]=8'b01101001;
   assign rom_data[4844]=8'b01101101;
   assign rom_data[4845]=8'b01100111;
   assign rom_data[4846]=8'b01101101;
   assign rom_data[4847]=8'b01100110;
   assign rom_data[4848]=8'b01101101;
   assign rom_data[4849]=8'b01100101;
   assign rom_data[4850]=8'b01101101;
   assign rom_data[4851]=8'b01100011;
   assign rom_data[4852]=8'b01101101;
   assign rom_data[4853]=8'b01100010;
   assign rom_data[4854]=8'b01101101;
   assign rom_data[4855]=8'b01100001;
   assign rom_data[4856]=8'b01101101;
   assign rom_data[4857]=8'b01011111;
   assign rom_data[4858]=8'b01101101;
   assign rom_data[4859]=8'b01011110;
   assign rom_data[4860]=8'b01101101;
   assign rom_data[4861]=8'b01011100;
   assign rom_data[4862]=8'b01101101;
   assign rom_data[4863]=8'b01011011;
   assign rom_data[4864]=8'b01101101;
   assign rom_data[4865]=8'b01011001;
   assign rom_data[4866]=8'b01101101;
   assign rom_data[4867]=8'b01011000;
   assign rom_data[4868]=8'b01101101;
   assign rom_data[4869]=8'b01010111;
   assign rom_data[4870]=8'b01101101;
   assign rom_data[4871]=8'b01010101;
   assign rom_data[4872]=8'b01101101;
   assign rom_data[4873]=8'b01010100;
   assign rom_data[4874]=8'b01101101;
   assign rom_data[4875]=8'b01010010;
   assign rom_data[4876]=8'b01101101;
   assign rom_data[4877]=8'b01010001;
   assign rom_data[4878]=8'b01101101;
   assign rom_data[4879]=8'b01010000;
   assign rom_data[4880]=8'b01101101;
   assign rom_data[4881]=8'b01001110;
   assign rom_data[4882]=8'b01101101;
   assign rom_data[4883]=8'b01001101;
   assign rom_data[4884]=8'b01101101;
   assign rom_data[4885]=8'b01001100;
   assign rom_data[4886]=8'b01101101;
   assign rom_data[4887]=8'b01001010;
   assign rom_data[4888]=8'b01101101;
   assign rom_data[4889]=8'b01001001;
   assign rom_data[4890]=8'b01101101;
   assign rom_data[4891]=8'b01001000;
   assign rom_data[4892]=8'b01101101;
   assign rom_data[4893]=8'b01000110;
   assign rom_data[4894]=8'b01101101;
   assign rom_data[4895]=8'b01000101;
   assign rom_data[4896]=8'b01101101;
   assign rom_data[4897]=8'b01000100;
   assign rom_data[4898]=8'b01101101;
   assign rom_data[4899]=8'b01000010;
   assign rom_data[4900]=8'b01101101;
   assign rom_data[4901]=8'b01000001;
   assign rom_data[4902]=8'b01101101;
   assign rom_data[4903]=8'b01000000;
   assign rom_data[4904]=8'b01101101;
   assign rom_data[4905]=8'b00111110;
   assign rom_data[4906]=8'b01101101;
   assign rom_data[4907]=8'b00111101;
   assign rom_data[4908]=8'b01101110;
   assign rom_data[4909]=8'b00111100;
   assign rom_data[4910]=8'b01101110;
   assign rom_data[4911]=8'b00111011;
   assign rom_data[4912]=8'b01101110;
   assign rom_data[4913]=8'b00111010;
   assign rom_data[4914]=8'b01101110;
   assign rom_data[4915]=8'b00111001;
   assign rom_data[4916]=8'b01101110;
   assign rom_data[4917]=8'b00111000;
   assign rom_data[4918]=8'b01101110;
   assign rom_data[4919]=8'b00110110;
   assign rom_data[4920]=8'b01101110;
   assign rom_data[4921]=8'b00110101;
   assign rom_data[4922]=8'b01101110;
   assign rom_data[4923]=8'b00110100;
   assign rom_data[4924]=8'b01101110;
   assign rom_data[4925]=8'b00110011;
   assign rom_data[4926]=8'b01101110;
   assign rom_data[4927]=8'b00110011;
   assign rom_data[4928]=8'b01101110;
   assign rom_data[4929]=8'b00110010;
   assign rom_data[4930]=8'b01101110;
   assign rom_data[4931]=8'b00110001;
   assign rom_data[4932]=8'b01101110;
   assign rom_data[4933]=8'b00110000;
   assign rom_data[4934]=8'b01101110;
   assign rom_data[4935]=8'b00101111;
   assign rom_data[4936]=8'b01101110;
   assign rom_data[4937]=8'b00101111;
   assign rom_data[4938]=8'b01101110;
   assign rom_data[4939]=8'b00101110;
   assign rom_data[4940]=8'b01101110;
   assign rom_data[4941]=8'b00101110;
   assign rom_data[4942]=8'b01101110;
   assign rom_data[4943]=8'b00101101;
   assign rom_data[4944]=8'b01101110;
   assign rom_data[4945]=8'b00101101;
   assign rom_data[4946]=8'b01101110;
   assign rom_data[4947]=8'b00101100;
   assign rom_data[4948]=8'b01101110;
   assign rom_data[4949]=8'b00101100;
   assign rom_data[4950]=8'b01101110;
   assign rom_data[4951]=8'b00101100;
   assign rom_data[4952]=8'b01101110;
   assign rom_data[4953]=8'b00101100;
   assign rom_data[4954]=8'b01101110;
   assign rom_data[4955]=8'b00101100;
   assign rom_data[4956]=8'b01101110;
   assign rom_data[4957]=8'b00101100;
   assign rom_data[4958]=8'b01101110;
   assign rom_data[4959]=8'b00101100;
   assign rom_data[4960]=8'b01101110;
   assign rom_data[4961]=8'b00101101;
   assign rom_data[4962]=8'b01101110;
   assign rom_data[4963]=8'b00101101;
   assign rom_data[4964]=8'b01101110;
   assign rom_data[4965]=8'b00101101;
   assign rom_data[4966]=8'b01101110;
   assign rom_data[4967]=8'b00101110;
   assign rom_data[4968]=8'b01101110;
   assign rom_data[4969]=8'b00101111;
   assign rom_data[4970]=8'b01101110;
   assign rom_data[4971]=8'b00101111;
   assign rom_data[4972]=8'b01101110;
   assign rom_data[4973]=8'b00110000;
   assign rom_data[4974]=8'b01101110;
   assign rom_data[4975]=8'b00110001;
   assign rom_data[4976]=8'b01101111;
   assign rom_data[4977]=8'b00110001;
   assign rom_data[4978]=8'b01101111;
   assign rom_data[4979]=8'b00110010;
   assign rom_data[4980]=8'b01101111;
   assign rom_data[4981]=8'b00110011;
   assign rom_data[4982]=8'b01101111;
   assign rom_data[4983]=8'b00110100;
   assign rom_data[4984]=8'b01101111;
   assign rom_data[4985]=8'b00110101;
   assign rom_data[4986]=8'b01101111;
   assign rom_data[4987]=8'b00110110;
   assign rom_data[4988]=8'b01101111;
   assign rom_data[4989]=8'b00110111;
   assign rom_data[4990]=8'b01101111;
   assign rom_data[4991]=8'b00111000;
   assign rom_data[4992]=8'b01101111;
   assign rom_data[4993]=8'b00111010;
   assign rom_data[4994]=8'b01101111;
   assign rom_data[4995]=8'b00111011;
   assign rom_data[4996]=8'b01101111;
   assign rom_data[4997]=8'b00111100;
   assign rom_data[4998]=8'b01101111;
   assign rom_data[4999]=8'b00111101;
   assign rom_data[5000]=8'b01101111;
   assign rom_data[5001]=8'b00111110;
   assign rom_data[5002]=8'b01101111;
   assign rom_data[5003]=8'b01000000;
   assign rom_data[5004]=8'b01101111;
   assign rom_data[5005]=8'b01000001;
   assign rom_data[5006]=8'b01101111;
   assign rom_data[5007]=8'b01000010;
   assign rom_data[5008]=8'b01101111;
   assign rom_data[5009]=8'b01000100;
   assign rom_data[5010]=8'b01101111;
   assign rom_data[5011]=8'b01000101;
   assign rom_data[5012]=8'b01101111;
   assign rom_data[5013]=8'b01000110;
   assign rom_data[5014]=8'b01101111;
   assign rom_data[5015]=8'b01001000;
   assign rom_data[5016]=8'b01101111;
   assign rom_data[5017]=8'b01001001;
   assign rom_data[5018]=8'b01101111;
   assign rom_data[5019]=8'b01001010;
   assign rom_data[5020]=8'b01101111;
   assign rom_data[5021]=8'b01001100;
   assign rom_data[5022]=8'b01101111;
   assign rom_data[5023]=8'b01001101;
   assign rom_data[5024]=8'b01101111;
   assign rom_data[5025]=8'b01001110;
   assign rom_data[5026]=8'b01101111;
   assign rom_data[5027]=8'b01010000;
   assign rom_data[5028]=8'b01101111;
   assign rom_data[5029]=8'b01010001;
   assign rom_data[5030]=8'b01101111;
   assign rom_data[5031]=8'b01010011;
   assign rom_data[5032]=8'b01101111;
   assign rom_data[5033]=8'b01010100;
   assign rom_data[5034]=8'b01101111;
   assign rom_data[5035]=8'b01010101;
   assign rom_data[5036]=8'b01101111;
   assign rom_data[5037]=8'b01010111;
   assign rom_data[5038]=8'b01101111;
   assign rom_data[5039]=8'b01011000;
   assign rom_data[5040]=8'b01101111;
   assign rom_data[5041]=8'b01011010;
   assign rom_data[5042]=8'b01101111;
   assign rom_data[5043]=8'b01011011;
   assign rom_data[5044]=8'b01101111;
   assign rom_data[5045]=8'b01011100;
   assign rom_data[5046]=8'b01101111;
   assign rom_data[5047]=8'b01011110;
   assign rom_data[5048]=8'b01101111;
   assign rom_data[5049]=8'b01011111;
   assign rom_data[5050]=8'b01101111;
   assign rom_data[5051]=8'b01100001;
   assign rom_data[5052]=8'b01101111;
   assign rom_data[5053]=8'b01100010;
   assign rom_data[5054]=8'b01101111;
   assign rom_data[5055]=8'b01100011;
   assign rom_data[5056]=8'b01110000;
   assign rom_data[5057]=8'b01100101;
   assign rom_data[5058]=8'b01110000;
   assign rom_data[5059]=8'b01100110;
   assign rom_data[5060]=8'b01110000;
   assign rom_data[5061]=8'b01101000;
   assign rom_data[5062]=8'b01110000;
   assign rom_data[5063]=8'b01101001;
   assign rom_data[5064]=8'b01110000;
   assign rom_data[5065]=8'b01101010;
   assign rom_data[5066]=8'b01110000;
   assign rom_data[5067]=8'b01101100;
   assign rom_data[5068]=8'b01110000;
   assign rom_data[5069]=8'b01101101;
   assign rom_data[5070]=8'b01110000;
   assign rom_data[5071]=8'b01101110;
   assign rom_data[5072]=8'b01110000;
   assign rom_data[5073]=8'b01110000;
   assign rom_data[5074]=8'b01110000;
   assign rom_data[5075]=8'b01110001;
   assign rom_data[5076]=8'b01110000;
   assign rom_data[5077]=8'b01110010;
   assign rom_data[5078]=8'b01110000;
   assign rom_data[5079]=8'b01110100;
   assign rom_data[5080]=8'b01110000;
   assign rom_data[5081]=8'b01110101;
   assign rom_data[5082]=8'b01110000;
   assign rom_data[5083]=8'b01110110;
   assign rom_data[5084]=8'b01110000;
   assign rom_data[5085]=8'b01110111;
   assign rom_data[5086]=8'b01110000;
   assign rom_data[5087]=8'b01111001;
   assign rom_data[5088]=8'b01110000;
   assign rom_data[5089]=8'b01111010;
   assign rom_data[5090]=8'b01110000;
   assign rom_data[5091]=8'b01111011;
   assign rom_data[5092]=8'b01110000;
   assign rom_data[5093]=8'b01111100;
   assign rom_data[5094]=8'b01110000;
   assign rom_data[5095]=8'b01111101;
   assign rom_data[5096]=8'b01110000;
   assign rom_data[5097]=8'b01111110;
   assign rom_data[5098]=8'b01110000;
   assign rom_data[5099]=8'b01111111;
   assign rom_data[5100]=8'b01110000;
   assign rom_data[5101]=8'b10000000;
   assign rom_data[5102]=8'b01110000;
   assign rom_data[5103]=8'b10000001;
   assign rom_data[5104]=8'b01110000;
   assign rom_data[5105]=8'b10000010;
   assign rom_data[5106]=8'b01110000;
   assign rom_data[5107]=8'b10000011;
   assign rom_data[5108]=8'b01110000;
   assign rom_data[5109]=8'b10000100;
   assign rom_data[5110]=8'b01110000;
   assign rom_data[5111]=8'b10000101;
   assign rom_data[5112]=8'b01110000;
   assign rom_data[5113]=8'b10000110;
   assign rom_data[5114]=8'b01110000;
   assign rom_data[5115]=8'b10000110;
   assign rom_data[5116]=8'b01110000;
   assign rom_data[5117]=8'b10000111;
   assign rom_data[5118]=8'b01110000;
   assign rom_data[5119]=8'b10001000;
   assign rom_data[5120]=8'b01110000;
   assign rom_data[5121]=8'b10001000;
   assign rom_data[5122]=8'b01110000;
   assign rom_data[5123]=8'b10001001;
   assign rom_data[5124]=8'b01110000;
   assign rom_data[5125]=8'b10001001;
   assign rom_data[5126]=8'b01110000;
   assign rom_data[5127]=8'b10001001;
   assign rom_data[5128]=8'b01110000;
   assign rom_data[5129]=8'b10001010;
   assign rom_data[5130]=8'b01110001;
   assign rom_data[5131]=8'b10001010;
   assign rom_data[5132]=8'b01110001;
   assign rom_data[5133]=8'b10001010;
   assign rom_data[5134]=8'b01110001;
   assign rom_data[5135]=8'b10001010;
   assign rom_data[5136]=8'b01110001;
   assign rom_data[5137]=8'b10001010;
   assign rom_data[5138]=8'b01110001;
   assign rom_data[5139]=8'b10001001;
   assign rom_data[5140]=8'b01110001;
   assign rom_data[5141]=8'b10001001;
   assign rom_data[5142]=8'b01110001;
   assign rom_data[5143]=8'b10001001;
   assign rom_data[5144]=8'b01110001;
   assign rom_data[5145]=8'b10001000;
   assign rom_data[5146]=8'b01110001;
   assign rom_data[5147]=8'b10001000;
   assign rom_data[5148]=8'b01110001;
   assign rom_data[5149]=8'b10000111;
   assign rom_data[5150]=8'b01110001;
   assign rom_data[5151]=8'b10000111;
   assign rom_data[5152]=8'b01110001;
   assign rom_data[5153]=8'b10000110;
   assign rom_data[5154]=8'b01110001;
   assign rom_data[5155]=8'b10000101;
   assign rom_data[5156]=8'b01110001;
   assign rom_data[5157]=8'b10000100;
   assign rom_data[5158]=8'b01110001;
   assign rom_data[5159]=8'b10000011;
   assign rom_data[5160]=8'b01110001;
   assign rom_data[5161]=8'b10000011;
   assign rom_data[5162]=8'b01110001;
   assign rom_data[5163]=8'b10000010;
   assign rom_data[5164]=8'b01110001;
   assign rom_data[5165]=8'b10000001;
   assign rom_data[5166]=8'b01110001;
   assign rom_data[5167]=8'b10000000;
   assign rom_data[5168]=8'b01110001;
   assign rom_data[5169]=8'b01111110;
   assign rom_data[5170]=8'b01110001;
   assign rom_data[5171]=8'b01111101;
   assign rom_data[5172]=8'b01110001;
   assign rom_data[5173]=8'b01111100;
   assign rom_data[5174]=8'b01110001;
   assign rom_data[5175]=8'b01111011;
   assign rom_data[5176]=8'b01110001;
   assign rom_data[5177]=8'b01111010;
   assign rom_data[5178]=8'b01110001;
   assign rom_data[5179]=8'b01111001;
   assign rom_data[5180]=8'b01110001;
   assign rom_data[5181]=8'b01110111;
   assign rom_data[5182]=8'b01110001;
   assign rom_data[5183]=8'b01110110;
   assign rom_data[5184]=8'b01110001;
   assign rom_data[5185]=8'b01110101;
   assign rom_data[5186]=8'b01110001;
   assign rom_data[5187]=8'b01110100;
   assign rom_data[5188]=8'b01110001;
   assign rom_data[5189]=8'b01110010;
   assign rom_data[5190]=8'b01110001;
   assign rom_data[5191]=8'b01110001;
   assign rom_data[5192]=8'b01110001;
   assign rom_data[5193]=8'b01110000;
   assign rom_data[5194]=8'b01110001;
   assign rom_data[5195]=8'b01101110;
   assign rom_data[5196]=8'b01110001;
   assign rom_data[5197]=8'b01101101;
   assign rom_data[5198]=8'b01110001;
   assign rom_data[5199]=8'b01101100;
   assign rom_data[5200]=8'b01110010;
   assign rom_data[5201]=8'b01101010;
   assign rom_data[5202]=8'b01110010;
   assign rom_data[5203]=8'b01101001;
   assign rom_data[5204]=8'b01110010;
   assign rom_data[5205]=8'b01100111;
   assign rom_data[5206]=8'b01110010;
   assign rom_data[5207]=8'b01100110;
   assign rom_data[5208]=8'b01110010;
   assign rom_data[5209]=8'b01100101;
   assign rom_data[5210]=8'b01110010;
   assign rom_data[5211]=8'b01100011;
   assign rom_data[5212]=8'b01110010;
   assign rom_data[5213]=8'b01100010;
   assign rom_data[5214]=8'b01110010;
   assign rom_data[5215]=8'b01100001;
   assign rom_data[5216]=8'b01110010;
   assign rom_data[5217]=8'b01011111;
   assign rom_data[5218]=8'b01110010;
   assign rom_data[5219]=8'b01011110;
   assign rom_data[5220]=8'b01110010;
   assign rom_data[5221]=8'b01011100;
   assign rom_data[5222]=8'b01110010;
   assign rom_data[5223]=8'b01011011;
   assign rom_data[5224]=8'b01110010;
   assign rom_data[5225]=8'b01011001;
   assign rom_data[5226]=8'b01110010;
   assign rom_data[5227]=8'b01011000;
   assign rom_data[5228]=8'b01110010;
   assign rom_data[5229]=8'b01010111;
   assign rom_data[5230]=8'b01110010;
   assign rom_data[5231]=8'b01010101;
   assign rom_data[5232]=8'b01110010;
   assign rom_data[5233]=8'b01010100;
   assign rom_data[5234]=8'b01110010;
   assign rom_data[5235]=8'b01010010;
   assign rom_data[5236]=8'b01110010;
   assign rom_data[5237]=8'b01010001;
   assign rom_data[5238]=8'b01110010;
   assign rom_data[5239]=8'b01010000;
   assign rom_data[5240]=8'b01110010;
   assign rom_data[5241]=8'b01001110;
   assign rom_data[5242]=8'b01110010;
   assign rom_data[5243]=8'b01001101;
   assign rom_data[5244]=8'b01110010;
   assign rom_data[5245]=8'b01001100;
   assign rom_data[5246]=8'b01110010;
   assign rom_data[5247]=8'b01001010;
   assign rom_data[5248]=8'b01110010;
   assign rom_data[5249]=8'b01001001;
   assign rom_data[5250]=8'b01110010;
   assign rom_data[5251]=8'b01001000;
   assign rom_data[5252]=8'b01110010;
   assign rom_data[5253]=8'b01000110;
   assign rom_data[5254]=8'b01110010;
   assign rom_data[5255]=8'b01000101;
   assign rom_data[5256]=8'b01110010;
   assign rom_data[5257]=8'b01000100;
   assign rom_data[5258]=8'b01110010;
   assign rom_data[5259]=8'b01000010;
   assign rom_data[5260]=8'b01110010;
   assign rom_data[5261]=8'b01000001;
   assign rom_data[5262]=8'b01110010;
   assign rom_data[5263]=8'b01000000;
   assign rom_data[5264]=8'b01110010;
   assign rom_data[5265]=8'b00111110;
   assign rom_data[5266]=8'b01110010;
   assign rom_data[5267]=8'b00111101;
   assign rom_data[5268]=8'b01110010;
   assign rom_data[5269]=8'b00111100;
   assign rom_data[5270]=8'b01110010;
   assign rom_data[5271]=8'b00111011;
   assign rom_data[5272]=8'b01110010;
   assign rom_data[5273]=8'b00111010;
   assign rom_data[5274]=8'b01110010;
   assign rom_data[5275]=8'b00111001;
   assign rom_data[5276]=8'b01110010;
   assign rom_data[5277]=8'b00111000;
   assign rom_data[5278]=8'b01110010;
   assign rom_data[5279]=8'b00110110;
   assign rom_data[5280]=8'b01110010;
   assign rom_data[5281]=8'b00110101;
   assign rom_data[5282]=8'b01110010;
   assign rom_data[5283]=8'b00110100;
   assign rom_data[5284]=8'b01110011;
   assign rom_data[5285]=8'b00110011;
   assign rom_data[5286]=8'b01110011;
   assign rom_data[5287]=8'b00110011;
   assign rom_data[5288]=8'b01110011;
   assign rom_data[5289]=8'b00110010;
   assign rom_data[5290]=8'b01110011;
   assign rom_data[5291]=8'b00110001;
   assign rom_data[5292]=8'b01110011;
   assign rom_data[5293]=8'b00110000;
   assign rom_data[5294]=8'b01110011;
   assign rom_data[5295]=8'b00101111;
   assign rom_data[5296]=8'b01110011;
   assign rom_data[5297]=8'b00101111;
   assign rom_data[5298]=8'b01110011;
   assign rom_data[5299]=8'b00101110;
   assign rom_data[5300]=8'b01110011;
   assign rom_data[5301]=8'b00101110;
   assign rom_data[5302]=8'b01110011;
   assign rom_data[5303]=8'b00101101;
   assign rom_data[5304]=8'b01110011;
   assign rom_data[5305]=8'b00101101;
   assign rom_data[5306]=8'b01110011;
   assign rom_data[5307]=8'b00101100;
   assign rom_data[5308]=8'b01110011;
   assign rom_data[5309]=8'b00101100;
   assign rom_data[5310]=8'b01110011;
   assign rom_data[5311]=8'b00101100;
   assign rom_data[5312]=8'b01110011;
   assign rom_data[5313]=8'b00101100;
   assign rom_data[5314]=8'b01110011;
   assign rom_data[5315]=8'b00101100;
   assign rom_data[5316]=8'b01110011;
   assign rom_data[5317]=8'b00101100;
   assign rom_data[5318]=8'b01110011;
   assign rom_data[5319]=8'b00101100;
   assign rom_data[5320]=8'b01110011;
   assign rom_data[5321]=8'b00101101;
   assign rom_data[5322]=8'b01110011;
   assign rom_data[5323]=8'b00101101;
   assign rom_data[5324]=8'b01110011;
   assign rom_data[5325]=8'b00101101;
   assign rom_data[5326]=8'b01110011;
   assign rom_data[5327]=8'b00101110;
   assign rom_data[5328]=8'b01110011;
   assign rom_data[5329]=8'b00101111;
   assign rom_data[5330]=8'b01110011;
   assign rom_data[5331]=8'b00101111;
   assign rom_data[5332]=8'b01110011;
   assign rom_data[5333]=8'b00110000;
   assign rom_data[5334]=8'b01110011;
   assign rom_data[5335]=8'b00110001;
   assign rom_data[5336]=8'b01110011;
   assign rom_data[5337]=8'b00110001;
   assign rom_data[5338]=8'b01110011;
   assign rom_data[5339]=8'b00110010;
   assign rom_data[5340]=8'b01110011;
   assign rom_data[5341]=8'b00110011;
   assign rom_data[5342]=8'b01110011;
   assign rom_data[5343]=8'b00110100;
   assign rom_data[5344]=8'b01110011;
   assign rom_data[5345]=8'b00110101;
   assign rom_data[5346]=8'b01110011;
   assign rom_data[5347]=8'b00110110;
   assign rom_data[5348]=8'b01110100;
   assign rom_data[5349]=8'b00110111;
   assign rom_data[5350]=8'b01110100;
   assign rom_data[5351]=8'b00111000;
   assign rom_data[5352]=8'b01110100;
   assign rom_data[5353]=8'b00111010;
   assign rom_data[5354]=8'b01110100;
   assign rom_data[5355]=8'b00111011;
   assign rom_data[5356]=8'b01110100;
   assign rom_data[5357]=8'b00111100;
   assign rom_data[5358]=8'b01110100;
   assign rom_data[5359]=8'b00111101;
   assign rom_data[5360]=8'b01110100;
   assign rom_data[5361]=8'b00111110;
   assign rom_data[5362]=8'b01110100;
   assign rom_data[5363]=8'b01000000;
   assign rom_data[5364]=8'b01110100;
   assign rom_data[5365]=8'b01000001;
   assign rom_data[5366]=8'b01110100;
   assign rom_data[5367]=8'b01000010;
   assign rom_data[5368]=8'b01110100;
   assign rom_data[5369]=8'b01000100;
   assign rom_data[5370]=8'b01110100;
   assign rom_data[5371]=8'b01000101;
   assign rom_data[5372]=8'b01110100;
   assign rom_data[5373]=8'b01000110;
   assign rom_data[5374]=8'b01110100;
   assign rom_data[5375]=8'b01001000;
   assign rom_data[5376]=8'b01110100;
   assign rom_data[5377]=8'b01001001;
   assign rom_data[5378]=8'b01110100;
   assign rom_data[5379]=8'b01001010;
   assign rom_data[5380]=8'b01110100;
   assign rom_data[5381]=8'b01001100;
   assign rom_data[5382]=8'b01110100;
   assign rom_data[5383]=8'b01001101;
   assign rom_data[5384]=8'b01110100;
   assign rom_data[5385]=8'b01001110;
   assign rom_data[5386]=8'b01110100;
   assign rom_data[5387]=8'b01010000;
   assign rom_data[5388]=8'b01110100;
   assign rom_data[5389]=8'b01010001;
   assign rom_data[5390]=8'b01110100;
   assign rom_data[5391]=8'b01010011;
   assign rom_data[5392]=8'b01110100;
   assign rom_data[5393]=8'b01010100;
   assign rom_data[5394]=8'b01110100;
   assign rom_data[5395]=8'b01010101;
   assign rom_data[5396]=8'b01110100;
   assign rom_data[5397]=8'b01010111;
   assign rom_data[5398]=8'b01110100;
   assign rom_data[5399]=8'b01011000;
   assign rom_data[5400]=8'b01110100;
   assign rom_data[5401]=8'b01011010;
   assign rom_data[5402]=8'b01110100;
   assign rom_data[5403]=8'b01011011;
   assign rom_data[5404]=8'b01110100;
   assign rom_data[5405]=8'b01011100;
   assign rom_data[5406]=8'b01110100;
   assign rom_data[5407]=8'b01011110;
   assign rom_data[5408]=8'b01110100;
   assign rom_data[5409]=8'b01011111;
   assign rom_data[5410]=8'b01110100;
   assign rom_data[5411]=8'b01100001;
   assign rom_data[5412]=8'b01110100;
   assign rom_data[5413]=8'b01100010;
   assign rom_data[5414]=8'b01110100;
   assign rom_data[5415]=8'b01100011;
   assign rom_data[5416]=8'b01110100;
   assign rom_data[5417]=8'b01100101;
   assign rom_data[5418]=8'b01110100;
   assign rom_data[5419]=8'b01100110;
   assign rom_data[5420]=8'b01110100;
   assign rom_data[5421]=8'b01101000;
   assign rom_data[5422]=8'b01110100;
   assign rom_data[5423]=8'b01101001;
   assign rom_data[5424]=8'b01110100;
   assign rom_data[5425]=8'b01101010;
   assign rom_data[5426]=8'b01110100;
   assign rom_data[5427]=8'b01101100;
   assign rom_data[5428]=8'b01110100;
   assign rom_data[5429]=8'b01101101;
   assign rom_data[5430]=8'b01110100;
   assign rom_data[5431]=8'b01101110;
   assign rom_data[5432]=8'b01110101;
   assign rom_data[5433]=8'b01110000;
   assign rom_data[5434]=8'b01110101;
   assign rom_data[5435]=8'b01110001;
   assign rom_data[5436]=8'b01110101;
   assign rom_data[5437]=8'b01110010;
   assign rom_data[5438]=8'b01110101;
   assign rom_data[5439]=8'b01110100;
   assign rom_data[5440]=8'b01110101;
   assign rom_data[5441]=8'b01110101;
   assign rom_data[5442]=8'b01110101;
   assign rom_data[5443]=8'b01110110;
   assign rom_data[5444]=8'b01110101;
   assign rom_data[5445]=8'b01110111;
   assign rom_data[5446]=8'b01110101;
   assign rom_data[5447]=8'b01111001;
   assign rom_data[5448]=8'b01110101;
   assign rom_data[5449]=8'b01111010;
   assign rom_data[5450]=8'b01110101;
   assign rom_data[5451]=8'b01111011;
   assign rom_data[5452]=8'b01110101;
   assign rom_data[5453]=8'b01111100;
   assign rom_data[5454]=8'b01110101;
   assign rom_data[5455]=8'b01111101;
   assign rom_data[5456]=8'b01110101;
   assign rom_data[5457]=8'b01111110;
   assign rom_data[5458]=8'b01110101;
   assign rom_data[5459]=8'b01111111;
   assign rom_data[5460]=8'b01110101;
   assign rom_data[5461]=8'b10000000;
   assign rom_data[5462]=8'b01110101;
   assign rom_data[5463]=8'b10000001;
   assign rom_data[5464]=8'b01110101;
   assign rom_data[5465]=8'b10000010;
   assign rom_data[5466]=8'b01110101;
   assign rom_data[5467]=8'b10000011;
   assign rom_data[5468]=8'b01110101;
   assign rom_data[5469]=8'b10000100;
   assign rom_data[5470]=8'b01110101;
   assign rom_data[5471]=8'b10000101;
   assign rom_data[5472]=8'b01110101;
   assign rom_data[5473]=8'b10000110;
   assign rom_data[5474]=8'b01110101;
   assign rom_data[5475]=8'b10000110;
   assign rom_data[5476]=8'b01110101;
   assign rom_data[5477]=8'b10000111;
   assign rom_data[5478]=8'b01110101;
   assign rom_data[5479]=8'b10001000;
   assign rom_data[5480]=8'b01110101;
   assign rom_data[5481]=8'b10001000;
   assign rom_data[5482]=8'b01110101;
   assign rom_data[5483]=8'b10001001;
   assign rom_data[5484]=8'b01110101;
   assign rom_data[5485]=8'b10001001;
   assign rom_data[5486]=8'b01110101;
   assign rom_data[5487]=8'b10001001;
   assign rom_data[5488]=8'b01110101;
   assign rom_data[5489]=8'b10001010;
   assign rom_data[5490]=8'b01110101;
   assign rom_data[5491]=8'b10001010;
   assign rom_data[5492]=8'b01110101;
   assign rom_data[5493]=8'b10001010;
   assign rom_data[5494]=8'b01110101;
   assign rom_data[5495]=8'b10001010;
   assign rom_data[5496]=8'b01110101;
   assign rom_data[5497]=8'b10001010;
   assign rom_data[5498]=8'b01110101;
   assign rom_data[5499]=8'b10001001;
   assign rom_data[5500]=8'b01110101;
   assign rom_data[5501]=8'b10001001;
   assign rom_data[5502]=8'b01110110;
   assign rom_data[5503]=8'b10001001;
   assign rom_data[5504]=8'b01110110;
   assign rom_data[5505]=8'b10001000;
   assign rom_data[5506]=8'b01110110;
   assign rom_data[5507]=8'b10001000;
   assign rom_data[5508]=8'b01110110;
   assign rom_data[5509]=8'b10000111;
   assign rom_data[5510]=8'b01110110;
   assign rom_data[5511]=8'b10000111;
   assign rom_data[5512]=8'b01110110;
   assign rom_data[5513]=8'b10000110;
   assign rom_data[5514]=8'b01110110;
   assign rom_data[5515]=8'b10000101;
   assign rom_data[5516]=8'b01110110;
   assign rom_data[5517]=8'b10000100;
   assign rom_data[5518]=8'b01110110;
   assign rom_data[5519]=8'b10000011;
   assign rom_data[5520]=8'b01110110;
   assign rom_data[5521]=8'b10000011;
   assign rom_data[5522]=8'b01110110;
   assign rom_data[5523]=8'b10000010;
   assign rom_data[5524]=8'b01110110;
   assign rom_data[5525]=8'b10000001;
   assign rom_data[5526]=8'b01110110;
   assign rom_data[5527]=8'b10000000;
   assign rom_data[5528]=8'b01110110;
   assign rom_data[5529]=8'b01111110;
   assign rom_data[5530]=8'b01110110;
   assign rom_data[5531]=8'b01111101;
   assign rom_data[5532]=8'b01110110;
   assign rom_data[5533]=8'b01111100;
   assign rom_data[5534]=8'b01110110;
   assign rom_data[5535]=8'b01111011;
   assign rom_data[5536]=8'b01110110;
   assign rom_data[5537]=8'b01111010;
   assign rom_data[5538]=8'b01110110;
   assign rom_data[5539]=8'b01111001;
   assign rom_data[5540]=8'b01110110;
   assign rom_data[5541]=8'b01110111;
   assign rom_data[5542]=8'b01110110;
   assign rom_data[5543]=8'b01110110;
   assign rom_data[5544]=8'b01110110;
   assign rom_data[5545]=8'b01110101;
   assign rom_data[5546]=8'b01110110;
   assign rom_data[5547]=8'b01110100;
   assign rom_data[5548]=8'b01110110;
   assign rom_data[5549]=8'b01110010;
   assign rom_data[5550]=8'b01110110;
   assign rom_data[5551]=8'b01110001;
   assign rom_data[5552]=8'b01110110;
   assign rom_data[5553]=8'b01110000;
   assign rom_data[5554]=8'b01110110;
   assign rom_data[5555]=8'b01101110;
   assign rom_data[5556]=8'b01110110;
   assign rom_data[5557]=8'b01101101;
   assign rom_data[5558]=8'b01110110;
   assign rom_data[5559]=8'b01101100;
   assign rom_data[5560]=8'b01110110;
   assign rom_data[5561]=8'b01101010;
   assign rom_data[5562]=8'b01110110;
   assign rom_data[5563]=8'b01101001;
   assign rom_data[5564]=8'b01110110;
   assign rom_data[5565]=8'b01100111;
   assign rom_data[5566]=8'b01110110;
   assign rom_data[5567]=8'b01100110;
   assign rom_data[5568]=8'b01110110;
   assign rom_data[5569]=8'b01100101;
   assign rom_data[5570]=8'b01110110;
   assign rom_data[5571]=8'b01100011;
   assign rom_data[5572]=8'b01110110;
   assign rom_data[5573]=8'b01100010;
   assign rom_data[5574]=8'b01110110;
   assign rom_data[5575]=8'b01100001;
   assign rom_data[5576]=8'b01110111;
   assign rom_data[5577]=8'b01011111;
   assign rom_data[5578]=8'b01110111;
   assign rom_data[5579]=8'b01011110;
   assign rom_data[5580]=8'b01110111;
   assign rom_data[5581]=8'b01011100;
   assign rom_data[5582]=8'b01110111;
   assign rom_data[5583]=8'b01011011;
   assign rom_data[5584]=8'b01110111;
   assign rom_data[5585]=8'b01011001;
   assign rom_data[5586]=8'b01110111;
   assign rom_data[5587]=8'b01011000;
   assign rom_data[5588]=8'b01110111;
   assign rom_data[5589]=8'b01010111;
   assign rom_data[5590]=8'b01110111;
   assign rom_data[5591]=8'b01010101;
   assign rom_data[5592]=8'b01110111;
   assign rom_data[5593]=8'b01010100;
   assign rom_data[5594]=8'b01110111;
   assign rom_data[5595]=8'b01010010;
   assign rom_data[5596]=8'b01110111;
   assign rom_data[5597]=8'b01010001;
   assign rom_data[5598]=8'b01110111;
   assign rom_data[5599]=8'b01010000;
   assign rom_data[5600]=8'b01110111;
   assign rom_data[5601]=8'b01001110;
   assign rom_data[5602]=8'b01110111;
   assign rom_data[5603]=8'b01001101;
   assign rom_data[5604]=8'b01110111;
   assign rom_data[5605]=8'b01001100;
   assign rom_data[5606]=8'b01110111;
   assign rom_data[5607]=8'b01001010;
   assign rom_data[5608]=8'b01110111;
   assign rom_data[5609]=8'b01001001;
   assign rom_data[5610]=8'b01110111;
   assign rom_data[5611]=8'b01001000;
   assign rom_data[5612]=8'b01110111;
   assign rom_data[5613]=8'b01000110;
   assign rom_data[5614]=8'b01110111;
   assign rom_data[5615]=8'b01000101;
   assign rom_data[5616]=8'b01110111;
   assign rom_data[5617]=8'b01000100;
   assign rom_data[5618]=8'b01110111;
   assign rom_data[5619]=8'b01000010;
   assign rom_data[5620]=8'b01110111;
   assign rom_data[5621]=8'b01000001;
   assign rom_data[5622]=8'b01110111;
   assign rom_data[5623]=8'b01000000;
   assign rom_data[5624]=8'b01110111;
   assign rom_data[5625]=8'b00111110;
   assign rom_data[5626]=8'b01110111;
   assign rom_data[5627]=8'b00111101;
   assign rom_data[5628]=8'b01110111;
   assign rom_data[5629]=8'b00111100;
   assign rom_data[5630]=8'b01110111;
   assign rom_data[5631]=8'b00111011;
   assign rom_data[5632]=8'b01110111;
   assign rom_data[5633]=8'b00111010;
   assign rom_data[5634]=8'b01110111;
   assign rom_data[5635]=8'b00111001;
   assign rom_data[5636]=8'b01110111;
   assign rom_data[5637]=8'b00111000;
   assign rom_data[5638]=8'b01110111;
   assign rom_data[5639]=8'b00110110;
   assign rom_data[5640]=8'b01110111;
   assign rom_data[5641]=8'b00110101;
   assign rom_data[5642]=8'b01110111;
   assign rom_data[5643]=8'b00110100;
   assign rom_data[5644]=8'b01110111;
   assign rom_data[5645]=8'b00110011;
   assign rom_data[5646]=8'b01110111;
   assign rom_data[5647]=8'b00110011;
   assign rom_data[5648]=8'b01110111;
   assign rom_data[5649]=8'b00110010;
   assign rom_data[5650]=8'b01110111;
   assign rom_data[5651]=8'b00110001;
   assign rom_data[5652]=8'b01110111;
   assign rom_data[5653]=8'b00110000;
   assign rom_data[5654]=8'b01110111;
   assign rom_data[5655]=8'b00101111;
   assign rom_data[5656]=8'b01111000;
   assign rom_data[5657]=8'b00101111;
   assign rom_data[5658]=8'b01111000;
   assign rom_data[5659]=8'b00101110;
   assign rom_data[5660]=8'b01111000;
   assign rom_data[5661]=8'b00101110;
   assign rom_data[5662]=8'b01111000;
   assign rom_data[5663]=8'b00101101;
   assign rom_data[5664]=8'b01111000;
   assign rom_data[5665]=8'b00101101;
   assign rom_data[5666]=8'b01111000;
   assign rom_data[5667]=8'b00101100;
   assign rom_data[5668]=8'b01111000;
   assign rom_data[5669]=8'b00101100;
   assign rom_data[5670]=8'b01111000;
   assign rom_data[5671]=8'b00101100;
   assign rom_data[5672]=8'b01111000;
   assign rom_data[5673]=8'b00101100;
   assign rom_data[5674]=8'b01111000;
   assign rom_data[5675]=8'b00101100;
   assign rom_data[5676]=8'b01111000;
   assign rom_data[5677]=8'b00101100;
   assign rom_data[5678]=8'b01111000;
   assign rom_data[5679]=8'b00101100;
   assign rom_data[5680]=8'b01111000;
   assign rom_data[5681]=8'b00101101;
   assign rom_data[5682]=8'b01111000;
   assign rom_data[5683]=8'b00101101;
   assign rom_data[5684]=8'b01111000;
   assign rom_data[5685]=8'b00101101;
   assign rom_data[5686]=8'b01111000;
   assign rom_data[5687]=8'b00101110;
   assign rom_data[5688]=8'b01111000;
   assign rom_data[5689]=8'b00101111;
   assign rom_data[5690]=8'b01111000;
   assign rom_data[5691]=8'b00101111;
   assign rom_data[5692]=8'b01111000;
   assign rom_data[5693]=8'b00110000;
   assign rom_data[5694]=8'b01111000;
   assign rom_data[5695]=8'b00110001;
   assign rom_data[5696]=8'b01111000;
   assign rom_data[5697]=8'b00110001;
   assign rom_data[5698]=8'b01111000;
   assign rom_data[5699]=8'b00110010;
   assign rom_data[5700]=8'b01111000;
   assign rom_data[5701]=8'b00110011;
   assign rom_data[5702]=8'b01111000;
   assign rom_data[5703]=8'b00110100;
   assign rom_data[5704]=8'b01111000;
   assign rom_data[5705]=8'b00110101;
   assign rom_data[5706]=8'b01111000;
   assign rom_data[5707]=8'b00110110;
   assign rom_data[5708]=8'b01111000;
   assign rom_data[5709]=8'b00110111;
   assign rom_data[5710]=8'b01111000;
   assign rom_data[5711]=8'b00111000;
   assign rom_data[5712]=8'b01111000;
   assign rom_data[5713]=8'b00111010;
   assign rom_data[5714]=8'b01111000;
   assign rom_data[5715]=8'b00111011;
   assign rom_data[5716]=8'b01111000;
   assign rom_data[5717]=8'b00111100;
   assign rom_data[5718]=8'b01111000;
   assign rom_data[5719]=8'b00111101;
   assign rom_data[5720]=8'b01111000;
   assign rom_data[5721]=8'b00111110;
   assign rom_data[5722]=8'b01111001;
   assign rom_data[5723]=8'b01000000;
   assign rom_data[5724]=8'b01111001;
   assign rom_data[5725]=8'b01000001;
   assign rom_data[5726]=8'b01111001;
   assign rom_data[5727]=8'b01000010;
   assign rom_data[5728]=8'b01111001;
   assign rom_data[5729]=8'b01000100;
   assign rom_data[5730]=8'b01111001;
   assign rom_data[5731]=8'b01000101;
   assign rom_data[5732]=8'b01111001;
   assign rom_data[5733]=8'b01000110;
   assign rom_data[5734]=8'b01111001;
   assign rom_data[5735]=8'b01001000;
   assign rom_data[5736]=8'b01111001;
   assign rom_data[5737]=8'b01001001;
   assign rom_data[5738]=8'b01111001;
   assign rom_data[5739]=8'b01001010;
   assign rom_data[5740]=8'b01111001;
   assign rom_data[5741]=8'b01001100;
   assign rom_data[5742]=8'b01111001;
   assign rom_data[5743]=8'b01001101;
   assign rom_data[5744]=8'b01111001;
   assign rom_data[5745]=8'b01001110;
   assign rom_data[5746]=8'b01111001;
   assign rom_data[5747]=8'b01010000;
   assign rom_data[5748]=8'b01111001;
   assign rom_data[5749]=8'b01010001;
   assign rom_data[5750]=8'b01111001;
   assign rom_data[5751]=8'b01010011;
   assign rom_data[5752]=8'b01111001;
   assign rom_data[5753]=8'b01010100;
   assign rom_data[5754]=8'b01111001;
   assign rom_data[5755]=8'b01010101;
   assign rom_data[5756]=8'b01111001;
   assign rom_data[5757]=8'b01010111;
   assign rom_data[5758]=8'b01111001;
   assign rom_data[5759]=8'b01011000;
   assign rom_data[5760]=8'b01111001;
   assign rom_data[5761]=8'b01011010;
   assign rom_data[5762]=8'b01111001;
   assign rom_data[5763]=8'b01011011;
   assign rom_data[5764]=8'b01111001;
   assign rom_data[5765]=8'b01011100;
   assign rom_data[5766]=8'b01111001;
   assign rom_data[5767]=8'b01011110;
   assign rom_data[5768]=8'b01111001;
   assign rom_data[5769]=8'b01011111;
   assign rom_data[5770]=8'b01111001;
   assign rom_data[5771]=8'b01100001;
   assign rom_data[5772]=8'b01111001;
   assign rom_data[5773]=8'b01100010;
   assign rom_data[5774]=8'b01111001;
   assign rom_data[5775]=8'b01100011;
   assign rom_data[5776]=8'b01111001;
   assign rom_data[5777]=8'b01100101;
   assign rom_data[5778]=8'b01111001;
   assign rom_data[5779]=8'b01100110;
   assign rom_data[5780]=8'b01111001;
   assign rom_data[5781]=8'b01101000;
   assign rom_data[5782]=8'b01111001;
   assign rom_data[5783]=8'b01101001;
   assign rom_data[5784]=8'b01111001;
   assign rom_data[5785]=8'b01101010;
   assign rom_data[5786]=8'b01111001;
   assign rom_data[5787]=8'b01101100;
   assign rom_data[5788]=8'b01111001;
   assign rom_data[5789]=8'b01101101;
   assign rom_data[5790]=8'b01111001;
   assign rom_data[5791]=8'b01101110;
   assign rom_data[5792]=8'b01111001;
   assign rom_data[5793]=8'b01110000;
   assign rom_data[5794]=8'b01111001;
   assign rom_data[5795]=8'b01110001;
   assign rom_data[5796]=8'b01111001;
   assign rom_data[5797]=8'b01110010;
   assign rom_data[5798]=8'b01111001;
   assign rom_data[5799]=8'b01110100;
   assign rom_data[5800]=8'b01111001;
   assign rom_data[5801]=8'b01110101;
   assign rom_data[5802]=8'b01111001;
   assign rom_data[5803]=8'b01110110;
   assign rom_data[5804]=8'b01111001;
   assign rom_data[5805]=8'b01110111;
   assign rom_data[5806]=8'b01111001;
   assign rom_data[5807]=8'b01111001;
   assign rom_data[5808]=8'b01111010;
   assign rom_data[5809]=8'b01111010;
   assign rom_data[5810]=8'b01111010;
   assign rom_data[5811]=8'b01111011;
   assign rom_data[5812]=8'b01111010;
   assign rom_data[5813]=8'b01111100;
   assign rom_data[5814]=8'b01111010;
   assign rom_data[5815]=8'b01111101;
   assign rom_data[5816]=8'b01111010;
   assign rom_data[5817]=8'b01111110;
   assign rom_data[5818]=8'b01111010;
   assign rom_data[5819]=8'b01111111;
   assign rom_data[5820]=8'b01111010;
   assign rom_data[5821]=8'b10000000;
   assign rom_data[5822]=8'b01111010;
   assign rom_data[5823]=8'b10000001;
   assign rom_data[5824]=8'b01111010;
   assign rom_data[5825]=8'b10000010;
   assign rom_data[5826]=8'b01111010;
   assign rom_data[5827]=8'b10000011;
   assign rom_data[5828]=8'b01111010;
   assign rom_data[5829]=8'b10000100;
   assign rom_data[5830]=8'b01111010;
   assign rom_data[5831]=8'b10000101;
   assign rom_data[5832]=8'b01111010;
   assign rom_data[5833]=8'b10000110;
   assign rom_data[5834]=8'b01111010;
   assign rom_data[5835]=8'b10000110;
   assign rom_data[5836]=8'b01111010;
   assign rom_data[5837]=8'b10000111;
   assign rom_data[5838]=8'b01111010;
   assign rom_data[5839]=8'b10001000;
   assign rom_data[5840]=8'b01111010;
   assign rom_data[5841]=8'b10001000;
   assign rom_data[5842]=8'b01111010;
   assign rom_data[5843]=8'b10001001;
   assign rom_data[5844]=8'b01111010;
   assign rom_data[5845]=8'b10001001;
   assign rom_data[5846]=8'b01111010;
   assign rom_data[5847]=8'b10001001;
   assign rom_data[5848]=8'b01111010;
   assign rom_data[5849]=8'b10001010;
   assign rom_data[5850]=8'b01111010;
   assign rom_data[5851]=8'b10001010;
   assign rom_data[5852]=8'b01111010;
   assign rom_data[5853]=8'b10001010;
   assign rom_data[5854]=8'b01111010;
   assign rom_data[5855]=8'b10001010;
   assign rom_data[5856]=8'b01111010;
   assign rom_data[5857]=8'b10001010;
   assign rom_data[5858]=8'b01111010;
   assign rom_data[5859]=8'b10001001;
   assign rom_data[5860]=8'b01111010;
   assign rom_data[5861]=8'b10001001;
   assign rom_data[5862]=8'b01111010;
   assign rom_data[5863]=8'b10001001;
   assign rom_data[5864]=8'b01111010;
   assign rom_data[5865]=8'b10001000;
   assign rom_data[5866]=8'b01111010;
   assign rom_data[5867]=8'b10001000;
   assign rom_data[5868]=8'b01111010;
   assign rom_data[5869]=8'b10000111;
   assign rom_data[5870]=8'b01111010;
   assign rom_data[5871]=8'b10000111;
   assign rom_data[5872]=8'b01111010;
   assign rom_data[5873]=8'b10000110;
   assign rom_data[5874]=8'b01111011;
   assign rom_data[5875]=8'b10000101;
   assign rom_data[5876]=8'b01111011;
   assign rom_data[5877]=8'b10000100;
   assign rom_data[5878]=8'b01111011;
   assign rom_data[5879]=8'b10000011;
   assign rom_data[5880]=8'b01111011;
   assign rom_data[5881]=8'b10000011;
   assign rom_data[5882]=8'b01111011;
   assign rom_data[5883]=8'b10000010;
   assign rom_data[5884]=8'b01111011;
   assign rom_data[5885]=8'b10000001;
   assign rom_data[5886]=8'b01111011;
   assign rom_data[5887]=8'b10000000;
   assign rom_data[5888]=8'b01111011;
   assign rom_data[5889]=8'b01111110;
   assign rom_data[5890]=8'b01111011;
   assign rom_data[5891]=8'b01111101;
   assign rom_data[5892]=8'b01111011;
   assign rom_data[5893]=8'b01111100;
   assign rom_data[5894]=8'b01111011;
   assign rom_data[5895]=8'b01111011;
   assign rom_data[5896]=8'b01111011;
   assign rom_data[5897]=8'b01111010;
   assign rom_data[5898]=8'b01111011;
   assign rom_data[5899]=8'b01111001;
   assign rom_data[5900]=8'b01111011;
   assign rom_data[5901]=8'b01110111;
   assign rom_data[5902]=8'b01111011;
   assign rom_data[5903]=8'b01110110;
   assign rom_data[5904]=8'b01111011;
   assign rom_data[5905]=8'b01110101;
   assign rom_data[5906]=8'b01111011;
   assign rom_data[5907]=8'b01110100;
   assign rom_data[5908]=8'b01111011;
   assign rom_data[5909]=8'b01110010;
   assign rom_data[5910]=8'b01111011;
   assign rom_data[5911]=8'b01110001;
   assign rom_data[5912]=8'b01111011;
   assign rom_data[5913]=8'b01110000;
   assign rom_data[5914]=8'b01111011;
   assign rom_data[5915]=8'b01101110;
   assign rom_data[5916]=8'b01111011;
   assign rom_data[5917]=8'b01101101;
   assign rom_data[5918]=8'b01111011;
   assign rom_data[5919]=8'b01101100;
   assign rom_data[5920]=8'b01111011;
   assign rom_data[5921]=8'b01101010;
   assign rom_data[5922]=8'b01111011;
   assign rom_data[5923]=8'b01101001;
   assign rom_data[5924]=8'b01111011;
   assign rom_data[5925]=8'b01100111;
   assign rom_data[5926]=8'b01111011;
   assign rom_data[5927]=8'b01100110;
   assign rom_data[5928]=8'b01111011;
   assign rom_data[5929]=8'b01100101;
   assign rom_data[5930]=8'b01111011;
   assign rom_data[5931]=8'b01100011;
   assign rom_data[5932]=8'b01111011;
   assign rom_data[5933]=8'b01100010;
   assign rom_data[5934]=8'b01111011;
   assign rom_data[5935]=8'b01100001;
   assign rom_data[5936]=8'b01111011;
   assign rom_data[5937]=8'b01011111;
   assign rom_data[5938]=8'b01111011;
   assign rom_data[5939]=8'b01011110;
   assign rom_data[5940]=8'b01111011;
   assign rom_data[5941]=8'b01011100;
   assign rom_data[5942]=8'b01111011;
   assign rom_data[5943]=8'b01011011;
   assign rom_data[5944]=8'b01111011;
   assign rom_data[5945]=8'b01011001;
   assign rom_data[5946]=8'b01111011;
   assign rom_data[5947]=8'b01011000;
   assign rom_data[5948]=8'b01111011;
   assign rom_data[5949]=8'b01010111;
   assign rom_data[5950]=8'b01111011;
   assign rom_data[5951]=8'b01010101;
   assign rom_data[5952]=8'b01111011;
   assign rom_data[5953]=8'b01010100;
   assign rom_data[5954]=8'b01111100;
   assign rom_data[5955]=8'b01010010;
   assign rom_data[5956]=8'b01111100;
   assign rom_data[5957]=8'b01010001;
   assign rom_data[5958]=8'b01111100;
   assign rom_data[5959]=8'b01010000;
   assign rom_data[5960]=8'b01111100;
   assign rom_data[5961]=8'b01001110;
   assign rom_data[5962]=8'b01111100;
   assign rom_data[5963]=8'b01001101;
   assign rom_data[5964]=8'b01111100;
   assign rom_data[5965]=8'b01001100;
   assign rom_data[5966]=8'b01111100;
   assign rom_data[5967]=8'b01001010;
   assign rom_data[5968]=8'b01111100;
   assign rom_data[5969]=8'b01001001;
   assign rom_data[5970]=8'b01111100;
   assign rom_data[5971]=8'b01001000;
   assign rom_data[5972]=8'b01111100;
   assign rom_data[5973]=8'b01000110;
   assign rom_data[5974]=8'b01111100;
   assign rom_data[5975]=8'b01000101;
   assign rom_data[5976]=8'b01111100;
   assign rom_data[5977]=8'b01000100;
   assign rom_data[5978]=8'b01111100;
   assign rom_data[5979]=8'b01000010;
   assign rom_data[5980]=8'b01111100;
   assign rom_data[5981]=8'b01000001;
   assign rom_data[5982]=8'b01111100;
   assign rom_data[5983]=8'b01000000;
   assign rom_data[5984]=8'b01111100;
   assign rom_data[5985]=8'b00111110;
   assign rom_data[5986]=8'b01111100;
   assign rom_data[5987]=8'b00111101;
   assign rom_data[5988]=8'b01111100;
   assign rom_data[5989]=8'b00111100;
   assign rom_data[5990]=8'b01111100;
   assign rom_data[5991]=8'b00111011;
   assign rom_data[5992]=8'b01111100;
   assign rom_data[5993]=8'b00111010;
   assign rom_data[5994]=8'b01111100;
   assign rom_data[5995]=8'b00111001;
   assign rom_data[5996]=8'b01111100;
   assign rom_data[5997]=8'b00111000;
   assign rom_data[5998]=8'b01111100;
   assign rom_data[5999]=8'b00110110;
   assign rom_data[6000]=8'b01111100;
   assign rom_data[6001]=8'b00110101;
   assign rom_data[6002]=8'b01111100;
   assign rom_data[6003]=8'b00110100;
   assign rom_data[6004]=8'b01111100;
   assign rom_data[6005]=8'b00110011;
   assign rom_data[6006]=8'b01111100;
   assign rom_data[6007]=8'b00110011;
   assign rom_data[6008]=8'b01111100;
   assign rom_data[6009]=8'b00110010;
   assign rom_data[6010]=8'b01111100;
   assign rom_data[6011]=8'b00110001;
   assign rom_data[6012]=8'b01111100;
   assign rom_data[6013]=8'b00110000;
   assign rom_data[6014]=8'b01111100;
   assign rom_data[6015]=8'b00101111;
   assign rom_data[6016]=8'b01111100;
   assign rom_data[6017]=8'b00101111;
   assign rom_data[6018]=8'b01111100;
   assign rom_data[6019]=8'b00101110;
   assign rom_data[6020]=8'b01111100;
   assign rom_data[6021]=8'b00101110;
   assign rom_data[6022]=8'b01111100;
   assign rom_data[6023]=8'b00101101;
   assign rom_data[6024]=8'b01111100;
   assign rom_data[6025]=8'b00101101;
   assign rom_data[6026]=8'b01111100;
   assign rom_data[6027]=8'b00101100;
   assign rom_data[6028]=8'b01111101;
   assign rom_data[6029]=8'b00101100;
   assign rom_data[6030]=8'b01111101;
   assign rom_data[6031]=8'b00101100;
   assign rom_data[6032]=8'b01111101;
   assign rom_data[6033]=8'b00101100;
   assign rom_data[6034]=8'b01111101;
   assign rom_data[6035]=8'b00101100;
   assign rom_data[6036]=8'b01111101;
   assign rom_data[6037]=8'b00101100;
   assign rom_data[6038]=8'b01111101;
   assign rom_data[6039]=8'b00101100;
   assign rom_data[6040]=8'b01111101;
   assign rom_data[6041]=8'b00101101;
   assign rom_data[6042]=8'b01111101;
   assign rom_data[6043]=8'b00101101;
   assign rom_data[6044]=8'b01111101;
   assign rom_data[6045]=8'b00101101;
   assign rom_data[6046]=8'b01111101;
   assign rom_data[6047]=8'b00101110;
   assign rom_data[6048]=8'b01111101;
   assign rom_data[6049]=8'b00101111;
   assign rom_data[6050]=8'b01111101;
   assign rom_data[6051]=8'b00101111;
   assign rom_data[6052]=8'b01111101;
   assign rom_data[6053]=8'b00110000;
   assign rom_data[6054]=8'b01111101;
   assign rom_data[6055]=8'b00110001;
   assign rom_data[6056]=8'b01111101;
   assign rom_data[6057]=8'b00110001;
   assign rom_data[6058]=8'b01111101;
   assign rom_data[6059]=8'b00110010;
   assign rom_data[6060]=8'b01111101;
   assign rom_data[6061]=8'b00110011;
   assign rom_data[6062]=8'b01111101;
   assign rom_data[6063]=8'b00110100;
   assign rom_data[6064]=8'b01111101;
   assign rom_data[6065]=8'b00110101;
   assign rom_data[6066]=8'b01111101;
   assign rom_data[6067]=8'b00110110;
   assign rom_data[6068]=8'b01111101;
   assign rom_data[6069]=8'b00110111;
   assign rom_data[6070]=8'b01111101;
   assign rom_data[6071]=8'b00111000;
   assign rom_data[6072]=8'b01111101;
   assign rom_data[6073]=8'b00111010;
   assign rom_data[6074]=8'b01111101;
   assign rom_data[6075]=8'b00111011;
   assign rom_data[6076]=8'b01111101;
   assign rom_data[6077]=8'b00111100;
   assign rom_data[6078]=8'b01111101;
   assign rom_data[6079]=8'b00111101;
   assign rom_data[6080]=8'b01111101;
   assign rom_data[6081]=8'b00111110;
   assign rom_data[6082]=8'b01111101;
   assign rom_data[6083]=8'b01000000;
   assign rom_data[6084]=8'b01111101;
   assign rom_data[6085]=8'b01000001;
   assign rom_data[6086]=8'b01111101;
   assign rom_data[6087]=8'b01000010;
   assign rom_data[6088]=8'b01111101;
   assign rom_data[6089]=8'b01000100;
   assign rom_data[6090]=8'b01111101;
   assign rom_data[6091]=8'b01000101;
   assign rom_data[6092]=8'b01111101;
   assign rom_data[6093]=8'b01000110;
   assign rom_data[6094]=8'b01111101;
   assign rom_data[6095]=8'b01001000;
   assign rom_data[6096]=8'b01111101;
   assign rom_data[6097]=8'b01001001;
   assign rom_data[6098]=8'b01111110;
   assign rom_data[6099]=8'b01001010;
   assign rom_data[6100]=8'b01111110;
   assign rom_data[6101]=8'b01001100;
   assign rom_data[6102]=8'b01111110;
   assign rom_data[6103]=8'b01001101;
   assign rom_data[6104]=8'b01111110;
   assign rom_data[6105]=8'b01001110;
   assign rom_data[6106]=8'b01111110;
   assign rom_data[6107]=8'b01010000;
   assign rom_data[6108]=8'b01111110;
   assign rom_data[6109]=8'b01010001;
   assign rom_data[6110]=8'b01111110;
   assign rom_data[6111]=8'b01010011;
   assign rom_data[6112]=8'b01111110;
   assign rom_data[6113]=8'b01010100;
   assign rom_data[6114]=8'b01111110;
   assign rom_data[6115]=8'b01010101;
   assign rom_data[6116]=8'b01111110;
   assign rom_data[6117]=8'b01010111;
   assign rom_data[6118]=8'b01111110;
   assign rom_data[6119]=8'b01011000;
   assign rom_data[6120]=8'b01111110;
   assign rom_data[6121]=8'b01011010;
   assign rom_data[6122]=8'b01111110;
   assign rom_data[6123]=8'b01011011;
   assign rom_data[6124]=8'b01111110;
   assign rom_data[6125]=8'b01011100;
   assign rom_data[6126]=8'b01111110;
   assign rom_data[6127]=8'b01011110;
   assign rom_data[6128]=8'b01111110;
   assign rom_data[6129]=8'b01011111;
   assign rom_data[6130]=8'b01111110;
   assign rom_data[6131]=8'b01100001;
   assign rom_data[6132]=8'b01111110;
   assign rom_data[6133]=8'b01100010;
   assign rom_data[6134]=8'b01111110;
   assign rom_data[6135]=8'b01100011;
   assign rom_data[6136]=8'b01111110;
   assign rom_data[6137]=8'b01100101;
   assign rom_data[6138]=8'b01111110;
   assign rom_data[6139]=8'b01100110;
   assign rom_data[6140]=8'b01111110;
   assign rom_data[6141]=8'b01101000;
   assign rom_data[6142]=8'b01111110;
   assign rom_data[6143]=8'b01101001;
   assign rom_data[6144]=8'b01111110;
   assign rom_data[6145]=8'b01101010;
   assign rom_data[6146]=8'b01111110;
   assign rom_data[6147]=8'b01101100;
   assign rom_data[6148]=8'b01111110;
   assign rom_data[6149]=8'b01101101;
   assign rom_data[6150]=8'b01111110;
   assign rom_data[6151]=8'b01101110;
   assign rom_data[6152]=8'b01111110;
   assign rom_data[6153]=8'b01110000;
   assign rom_data[6154]=8'b01111110;
   assign rom_data[6155]=8'b01110001;
   assign rom_data[6156]=8'b01111110;
   assign rom_data[6157]=8'b01110010;
   assign rom_data[6158]=8'b01111110;
   assign rom_data[6159]=8'b01110100;
   assign rom_data[6160]=8'b01111110;
   assign rom_data[6161]=8'b01110101;
   assign rom_data[6162]=8'b01111110;
   assign rom_data[6163]=8'b01110110;
   assign rom_data[6164]=8'b01111110;
   assign rom_data[6165]=8'b01110111;
   assign rom_data[6166]=8'b01111110;
   assign rom_data[6167]=8'b01111001;
   assign rom_data[6168]=8'b01111110;
   assign rom_data[6169]=8'b01111010;
   assign rom_data[6170]=8'b01111110;
   assign rom_data[6171]=8'b01111011;
   assign rom_data[6172]=8'b01111110;
   assign rom_data[6173]=8'b01111100;
   assign rom_data[6174]=8'b01111110;
   assign rom_data[6175]=8'b01111101;
   assign rom_data[6176]=8'b01111110;
   assign rom_data[6177]=8'b01111110;
   assign rom_data[6178]=8'b01111110;
   assign rom_data[6179]=8'b01111111;
   assign rom_data[6180]=8'b01111110;
   assign rom_data[6181]=8'b10000000;
   assign rom_data[6182]=8'b01111111;
   assign rom_data[6183]=8'b10000001;
   assign rom_data[6184]=8'b01111111;
   assign rom_data[6185]=8'b10000010;
   assign rom_data[6186]=8'b01111111;
   assign rom_data[6187]=8'b10000011;
   assign rom_data[6188]=8'b01111111;
   assign rom_data[6189]=8'b10000100;
   assign rom_data[6190]=8'b01111111;
   assign rom_data[6191]=8'b10000101;
   assign rom_data[6192]=8'b01111111;
   assign rom_data[6193]=8'b10000110;
   assign rom_data[6194]=8'b01111111;
   assign rom_data[6195]=8'b10000110;
   assign rom_data[6196]=8'b01111111;
   assign rom_data[6197]=8'b10000111;
   assign rom_data[6198]=8'b01111111;
   assign rom_data[6199]=8'b10001000;
   assign rom_data[6200]=8'b01111111;
   assign rom_data[6201]=8'b10001000;
   assign rom_data[6202]=8'b01111111;
   assign rom_data[6203]=8'b10001001;
   assign rom_data[6204]=8'b01111111;
   assign rom_data[6205]=8'b10001001;
   assign rom_data[6206]=8'b01111111;
   assign rom_data[6207]=8'b10001001;
   assign rom_data[6208]=8'b01111111;
   assign rom_data[6209]=8'b10001010;
   assign rom_data[6210]=8'b01111111;
   assign rom_data[6211]=8'b10001010;
   assign rom_data[6212]=8'b01111111;
   assign rom_data[6213]=8'b10001010;
   assign rom_data[6214]=8'b01111111;
   assign rom_data[6215]=8'b10001010;
   assign rom_data[6216]=8'b01111111;
   assign rom_data[6217]=8'b10001010;
   assign rom_data[6218]=8'b01111111;
   assign rom_data[6219]=8'b10001001;
   assign rom_data[6220]=8'b01111111;
   assign rom_data[6221]=8'b10001001;
   assign rom_data[6222]=8'b01111111;
   assign rom_data[6223]=8'b10001001;
   assign rom_data[6224]=8'b01111111;
   assign rom_data[6225]=8'b10001000;
   assign rom_data[6226]=8'b01111111;
   assign rom_data[6227]=8'b10001000;
   assign rom_data[6228]=8'b01111111;
   assign rom_data[6229]=8'b10000111;
   assign rom_data[6230]=8'b01111111;
   assign rom_data[6231]=8'b10000111;
   assign rom_data[6232]=8'b01111111;
   assign rom_data[6233]=8'b10000110;
   assign rom_data[6234]=8'b01111111;
   assign rom_data[6235]=8'b10000101;
   assign rom_data[6236]=8'b01111111;
   assign rom_data[6237]=8'b10000100;
   assign rom_data[6238]=8'b01111111;
   assign rom_data[6239]=8'b10000011;
   assign rom_data[6240]=8'b01111111;
   assign rom_data[6241]=8'b10000011;
   assign rom_data[6242]=8'b01111111;
   assign rom_data[6243]=8'b10000010;
   assign rom_data[6244]=8'b01111111;
   assign rom_data[6245]=8'b10000001;
   assign rom_data[6246]=8'b10000000;
   assign rom_data[6247]=8'b10000000;
   assign rom_data[6248]=8'b10000000;
   assign rom_data[6249]=8'b01111110;
   assign rom_data[6250]=8'b10000000;
   assign rom_data[6251]=8'b01111101;
   assign rom_data[6252]=8'b10000000;
   assign rom_data[6253]=8'b01111100;
   assign rom_data[6254]=8'b10000000;
   assign rom_data[6255]=8'b01111011;
   assign rom_data[6256]=8'b10000000;
   assign rom_data[6257]=8'b01111010;
   assign rom_data[6258]=8'b10000000;
   assign rom_data[6259]=8'b01111001;
   assign rom_data[6260]=8'b10000000;
   assign rom_data[6261]=8'b01110111;
   assign rom_data[6262]=8'b10000000;
   assign rom_data[6263]=8'b01110110;
   assign rom_data[6264]=8'b10000000;
   assign rom_data[6265]=8'b01110101;
   assign rom_data[6266]=8'b10000000;
   assign rom_data[6267]=8'b01110100;
   assign rom_data[6268]=8'b10000000;
   assign rom_data[6269]=8'b01110010;
   assign rom_data[6270]=8'b10000000;
   assign rom_data[6271]=8'b01110001;
   assign rom_data[6272]=8'b10000000;
   assign rom_data[6273]=8'b01110000;
   assign rom_data[6274]=8'b10000000;
   assign rom_data[6275]=8'b01101110;
   assign rom_data[6276]=8'b10000000;
   assign rom_data[6277]=8'b01101101;
   assign rom_data[6278]=8'b10000000;
   assign rom_data[6279]=8'b01101100;
   assign rom_data[6280]=8'b10000000;
   assign rom_data[6281]=8'b01101010;
   assign rom_data[6282]=8'b10000000;
   assign rom_data[6283]=8'b01101001;
   assign rom_data[6284]=8'b10000000;
   assign rom_data[6285]=8'b01100111;
   assign rom_data[6286]=8'b10000000;
   assign rom_data[6287]=8'b01100110;
   assign rom_data[6288]=8'b10000000;
   assign rom_data[6289]=8'b01100101;
   assign rom_data[6290]=8'b10000000;
   assign rom_data[6291]=8'b01100011;
   assign rom_data[6292]=8'b10000000;
   assign rom_data[6293]=8'b01100010;
   assign rom_data[6294]=8'b10000000;
   assign rom_data[6295]=8'b01100001;
   assign rom_data[6296]=8'b10000000;
   assign rom_data[6297]=8'b01011111;
   assign rom_data[6298]=8'b10000000;
   assign rom_data[6299]=8'b01011110;
   assign rom_data[6300]=8'b10000000;
   assign rom_data[6301]=8'b01011100;
   assign rom_data[6302]=8'b10000000;
   assign rom_data[6303]=8'b01011011;
   assign rom_data[6304]=8'b10000000;
   assign rom_data[6305]=8'b01011001;
   assign rom_data[6306]=8'b10000000;
   assign rom_data[6307]=8'b01011000;
   assign rom_data[6308]=8'b10000000;
   assign rom_data[6309]=8'b01010111;
   assign rom_data[6310]=8'b10000000;
   assign rom_data[6311]=8'b01010101;
   assign rom_data[6312]=8'b10000000;
   assign rom_data[6313]=8'b01010100;
   assign rom_data[6314]=8'b10000000;
   assign rom_data[6315]=8'b01010010;
   assign rom_data[6316]=8'b10000000;
   assign rom_data[6317]=8'b01010001;
   assign rom_data[6318]=8'b10000000;
   assign rom_data[6319]=8'b01010000;
   assign rom_data[6320]=8'b10000000;
   assign rom_data[6321]=8'b01001110;
   assign rom_data[6322]=8'b10000000;
   assign rom_data[6323]=8'b01001101;
   assign rom_data[6324]=8'b10000000;
   assign rom_data[6325]=8'b01001100;
   assign rom_data[6326]=8'b10000000;
   assign rom_data[6327]=8'b01001010;
   assign rom_data[6328]=8'b10000000;
   assign rom_data[6329]=8'b01001001;
   assign rom_data[6330]=8'b10000001;
   assign rom_data[6331]=8'b01001000;
   assign rom_data[6332]=8'b10000001;
   assign rom_data[6333]=8'b01000110;
   assign rom_data[6334]=8'b10000001;
   assign rom_data[6335]=8'b01000101;
   assign rom_data[6336]=8'b10000001;
   assign rom_data[6337]=8'b01000100;
   assign rom_data[6338]=8'b10000001;
   assign rom_data[6339]=8'b01000010;
   assign rom_data[6340]=8'b10000001;
   assign rom_data[6341]=8'b01000001;
   assign rom_data[6342]=8'b10000001;
   assign rom_data[6343]=8'b01000000;
   assign rom_data[6344]=8'b10000001;
   assign rom_data[6345]=8'b00111110;
   assign rom_data[6346]=8'b10000001;
   assign rom_data[6347]=8'b00111101;
   assign rom_data[6348]=8'b10000001;
   assign rom_data[6349]=8'b00111100;
   assign rom_data[6350]=8'b10000001;
   assign rom_data[6351]=8'b00111011;
   assign rom_data[6352]=8'b10000001;
   assign rom_data[6353]=8'b00111010;
   assign rom_data[6354]=8'b10000001;
   assign rom_data[6355]=8'b00111001;
   assign rom_data[6356]=8'b10000001;
   assign rom_data[6357]=8'b00111000;
   assign rom_data[6358]=8'b10000001;
   assign rom_data[6359]=8'b00110110;
   assign rom_data[6360]=8'b10000001;
   assign rom_data[6361]=8'b00110101;
   assign rom_data[6362]=8'b10000001;
   assign rom_data[6363]=8'b00110100;
   assign rom_data[6364]=8'b10000001;
   assign rom_data[6365]=8'b00110011;
   assign rom_data[6366]=8'b10000001;
   assign rom_data[6367]=8'b00110011;
   assign rom_data[6368]=8'b10000001;
   assign rom_data[6369]=8'b00110010;
   assign rom_data[6370]=8'b10000001;
   assign rom_data[6371]=8'b00110001;
   assign rom_data[6372]=8'b10000001;
   assign rom_data[6373]=8'b00110000;
   assign rom_data[6374]=8'b10000001;
   assign rom_data[6375]=8'b00101111;
   assign rom_data[6376]=8'b10000001;
   assign rom_data[6377]=8'b00101111;
   assign rom_data[6378]=8'b10000001;
   assign rom_data[6379]=8'b00101110;
   assign rom_data[6380]=8'b10000001;
   assign rom_data[6381]=8'b00101110;
   assign rom_data[6382]=8'b10000001;
   assign rom_data[6383]=8'b00101101;
   assign rom_data[6384]=8'b10000001;
   assign rom_data[6385]=8'b00101101;
   assign rom_data[6386]=8'b10000001;
   assign rom_data[6387]=8'b00101100;
   assign rom_data[6388]=8'b10000001;
   assign rom_data[6389]=8'b00101100;
   assign rom_data[6390]=8'b10000001;
   assign rom_data[6391]=8'b00101100;
   assign rom_data[6392]=8'b10000001;
   assign rom_data[6393]=8'b00101100;
   assign rom_data[6394]=8'b10000001;
   assign rom_data[6395]=8'b00101100;
   assign rom_data[6396]=8'b10000001;
   assign rom_data[6397]=8'b00101100;
   assign rom_data[6398]=8'b10000001;
   assign rom_data[6399]=8'b00101100;
   assign rom_data[6400]=8'b10000010;
   assign rom_data[6401]=8'b00101101;
   assign rom_data[6402]=8'b10000010;
   assign rom_data[6403]=8'b00101101;
   assign rom_data[6404]=8'b10000010;
   assign rom_data[6405]=8'b00101101;
   assign rom_data[6406]=8'b10000010;
   assign rom_data[6407]=8'b00101110;
   assign rom_data[6408]=8'b10000010;
   assign rom_data[6409]=8'b00101111;
   assign rom_data[6410]=8'b10000010;
   assign rom_data[6411]=8'b00101111;
   assign rom_data[6412]=8'b10000010;
   assign rom_data[6413]=8'b00110000;
   assign rom_data[6414]=8'b10000010;
   assign rom_data[6415]=8'b00110001;
   assign rom_data[6416]=8'b10000010;
   assign rom_data[6417]=8'b00110001;
   assign rom_data[6418]=8'b10000010;
   assign rom_data[6419]=8'b00110010;
   assign rom_data[6420]=8'b10000010;
   assign rom_data[6421]=8'b00110011;
   assign rom_data[6422]=8'b10000010;
   assign rom_data[6423]=8'b00110100;
   assign rom_data[6424]=8'b10000010;
   assign rom_data[6425]=8'b00110101;
   assign rom_data[6426]=8'b10000010;
   assign rom_data[6427]=8'b00110110;
   assign rom_data[6428]=8'b10000010;
   assign rom_data[6429]=8'b00110111;
   assign rom_data[6430]=8'b10000010;
   assign rom_data[6431]=8'b00111000;
   assign rom_data[6432]=8'b10000010;
   assign rom_data[6433]=8'b00111010;
   assign rom_data[6434]=8'b10000010;
   assign rom_data[6435]=8'b00111011;
   assign rom_data[6436]=8'b10000010;
   assign rom_data[6437]=8'b00111100;
   assign rom_data[6438]=8'b10000010;
   assign rom_data[6439]=8'b00111101;
   assign rom_data[6440]=8'b10000010;
   assign rom_data[6441]=8'b00111110;
   assign rom_data[6442]=8'b10000010;
   assign rom_data[6443]=8'b01000000;
   assign rom_data[6444]=8'b10000010;
   assign rom_data[6445]=8'b01000001;
   assign rom_data[6446]=8'b10000010;
   assign rom_data[6447]=8'b01000010;
   assign rom_data[6448]=8'b10000010;
   assign rom_data[6449]=8'b01000100;
   assign rom_data[6450]=8'b10000010;
   assign rom_data[6451]=8'b01000101;
   assign rom_data[6452]=8'b10000010;
   assign rom_data[6453]=8'b01000110;
   assign rom_data[6454]=8'b10000010;
   assign rom_data[6455]=8'b01001000;
   assign rom_data[6456]=8'b10000010;
   assign rom_data[6457]=8'b01001001;
   assign rom_data[6458]=8'b10000010;
   assign rom_data[6459]=8'b01001010;
   assign rom_data[6460]=8'b10000010;
   assign rom_data[6461]=8'b01001100;
   assign rom_data[6462]=8'b10000010;
   assign rom_data[6463]=8'b01001101;
   assign rom_data[6464]=8'b10000010;
   assign rom_data[6465]=8'b01001110;
   assign rom_data[6466]=8'b10000010;
   assign rom_data[6467]=8'b01010000;
   assign rom_data[6468]=8'b10000010;
   assign rom_data[6469]=8'b01010001;
   assign rom_data[6470]=8'b10000010;
   assign rom_data[6471]=8'b01010011;
   assign rom_data[6472]=8'b10000010;
   assign rom_data[6473]=8'b01010100;
   assign rom_data[6474]=8'b10000011;
   assign rom_data[6475]=8'b01010101;
   assign rom_data[6476]=8'b10000011;
   assign rom_data[6477]=8'b01010111;
   assign rom_data[6478]=8'b10000011;
   assign rom_data[6479]=8'b01011000;
   assign rom_data[6480]=8'b10000011;
   assign rom_data[6481]=8'b01011010;
   assign rom_data[6482]=8'b10000011;
   assign rom_data[6483]=8'b01011011;
   assign rom_data[6484]=8'b10000011;
   assign rom_data[6485]=8'b01011100;
   assign rom_data[6486]=8'b10000011;
   assign rom_data[6487]=8'b01011110;
   assign rom_data[6488]=8'b10000011;
   assign rom_data[6489]=8'b01011111;
   assign rom_data[6490]=8'b10000011;
   assign rom_data[6491]=8'b01100001;
   assign rom_data[6492]=8'b10000011;
   assign rom_data[6493]=8'b01100010;
   assign rom_data[6494]=8'b10000011;
   assign rom_data[6495]=8'b01100011;
   assign rom_data[6496]=8'b10000011;
   assign rom_data[6497]=8'b01100101;
   assign rom_data[6498]=8'b10000011;
   assign rom_data[6499]=8'b01100110;
   assign rom_data[6500]=8'b10000011;
   assign rom_data[6501]=8'b01101000;
   assign rom_data[6502]=8'b10000011;
   assign rom_data[6503]=8'b01101001;
   assign rom_data[6504]=8'b10000011;
   assign rom_data[6505]=8'b01101010;
   assign rom_data[6506]=8'b10000011;
   assign rom_data[6507]=8'b01101100;
   assign rom_data[6508]=8'b10000011;
   assign rom_data[6509]=8'b01101101;
   assign rom_data[6510]=8'b10000011;
   assign rom_data[6511]=8'b01101110;
   assign rom_data[6512]=8'b10000011;
   assign rom_data[6513]=8'b01110000;
   assign rom_data[6514]=8'b10000011;
   assign rom_data[6515]=8'b01110001;
   assign rom_data[6516]=8'b10000011;
   assign rom_data[6517]=8'b01110010;
   assign rom_data[6518]=8'b10000011;
   assign rom_data[6519]=8'b01110100;
   assign rom_data[6520]=8'b10000011;
   assign rom_data[6521]=8'b01110101;
   assign rom_data[6522]=8'b10000011;
   assign rom_data[6523]=8'b01110110;
   assign rom_data[6524]=8'b10000011;
   assign rom_data[6525]=8'b01110111;
   assign rom_data[6526]=8'b10000011;
   assign rom_data[6527]=8'b01111001;
   assign rom_data[6528]=8'b10000011;
   assign rom_data[6529]=8'b01111010;
   assign rom_data[6530]=8'b10000011;
   assign rom_data[6531]=8'b01111011;
   assign rom_data[6532]=8'b10000011;
   assign rom_data[6533]=8'b01111100;
   assign rom_data[6534]=8'b10000011;
   assign rom_data[6535]=8'b01111101;
   assign rom_data[6536]=8'b10000011;
   assign rom_data[6537]=8'b01111110;
   assign rom_data[6538]=8'b10000011;
   assign rom_data[6539]=8'b01111111;
   assign rom_data[6540]=8'b10000011;
   assign rom_data[6541]=8'b10000000;
   assign rom_data[6542]=8'b10000011;
   assign rom_data[6543]=8'b10000001;
   assign rom_data[6544]=8'b10000011;
   assign rom_data[6545]=8'b10000010;
   assign rom_data[6546]=8'b10000011;
   assign rom_data[6547]=8'b10000011;
   assign rom_data[6548]=8'b10000011;
   assign rom_data[6549]=8'b10000100;
   assign rom_data[6550]=8'b10000011;
   assign rom_data[6551]=8'b10000101;
   assign rom_data[6552]=8'b10000011;
   assign rom_data[6553]=8'b10000110;
   assign rom_data[6554]=8'b10000100;
   assign rom_data[6555]=8'b10000110;
   assign rom_data[6556]=8'b10000100;
   assign rom_data[6557]=8'b10000111;
   assign rom_data[6558]=8'b10000100;
   assign rom_data[6559]=8'b10001000;
   assign rom_data[6560]=8'b10000100;
   assign rom_data[6561]=8'b10001000;
   assign rom_data[6562]=8'b10000100;
   assign rom_data[6563]=8'b10001001;
   assign rom_data[6564]=8'b10000100;
   assign rom_data[6565]=8'b10001001;
   assign rom_data[6566]=8'b10000100;
   assign rom_data[6567]=8'b10001001;
   assign rom_data[6568]=8'b10000100;
   assign rom_data[6569]=8'b10001010;
   assign rom_data[6570]=8'b10000100;
   assign rom_data[6571]=8'b10001010;
   assign rom_data[6572]=8'b10000100;
   assign rom_data[6573]=8'b10001010;
   assign rom_data[6574]=8'b10000100;
   assign rom_data[6575]=8'b10001010;
   assign rom_data[6576]=8'b10000100;
   assign rom_data[6577]=8'b10001010;
   assign rom_data[6578]=8'b10000100;
   assign rom_data[6579]=8'b10001001;
   assign rom_data[6580]=8'b10000100;
   assign rom_data[6581]=8'b10001001;
   assign rom_data[6582]=8'b10000100;
   assign rom_data[6583]=8'b10001001;
   assign rom_data[6584]=8'b10000100;
   assign rom_data[6585]=8'b10001000;
   assign rom_data[6586]=8'b10000100;
   assign rom_data[6587]=8'b10001000;
   assign rom_data[6588]=8'b10000100;
   assign rom_data[6589]=8'b10000111;
   assign rom_data[6590]=8'b10000100;
   assign rom_data[6591]=8'b10000111;
   assign rom_data[6592]=8'b10000100;
   assign rom_data[6593]=8'b10000110;
   assign rom_data[6594]=8'b10000100;
   assign rom_data[6595]=8'b10000101;
   assign rom_data[6596]=8'b10000100;
   assign rom_data[6597]=8'b10000100;
   assign rom_data[6598]=8'b10000100;
   assign rom_data[6599]=8'b10000011;
   assign rom_data[6600]=8'b10000100;
   assign rom_data[6601]=8'b10000011;
   assign rom_data[6602]=8'b10000100;
   assign rom_data[6603]=8'b10000010;
   assign rom_data[6604]=8'b10000100;
   assign rom_data[6605]=8'b10000001;
   assign rom_data[6606]=8'b10000100;
   assign rom_data[6607]=8'b10000000;
   assign rom_data[6608]=8'b10000100;
   assign rom_data[6609]=8'b01111110;
   assign rom_data[6610]=8'b10000100;
   assign rom_data[6611]=8'b01111101;
   assign rom_data[6612]=8'b10000100;
   assign rom_data[6613]=8'b01111100;
   assign rom_data[6614]=8'b10000100;
   assign rom_data[6615]=8'b01111011;
   assign rom_data[6616]=8'b10000100;
   assign rom_data[6617]=8'b01111010;
   assign rom_data[6618]=8'b10000100;
   assign rom_data[6619]=8'b01111001;
   assign rom_data[6620]=8'b10000100;
   assign rom_data[6621]=8'b01110111;
   assign rom_data[6622]=8'b10000101;
   assign rom_data[6623]=8'b01110110;
   assign rom_data[6624]=8'b10000101;
   assign rom_data[6625]=8'b01110101;
   assign rom_data[6626]=8'b10000101;
   assign rom_data[6627]=8'b01110100;
   assign rom_data[6628]=8'b10000101;
   assign rom_data[6629]=8'b01110010;
   assign rom_data[6630]=8'b10000101;
   assign rom_data[6631]=8'b01110001;
   assign rom_data[6632]=8'b10000101;
   assign rom_data[6633]=8'b01110000;
   assign rom_data[6634]=8'b10000101;
   assign rom_data[6635]=8'b01101110;
   assign rom_data[6636]=8'b10000101;
   assign rom_data[6637]=8'b01101101;
   assign rom_data[6638]=8'b10000101;
   assign rom_data[6639]=8'b01101100;
   assign rom_data[6640]=8'b10000101;
   assign rom_data[6641]=8'b01101010;
   assign rom_data[6642]=8'b10000101;
   assign rom_data[6643]=8'b01101001;
   assign rom_data[6644]=8'b10000101;
   assign rom_data[6645]=8'b01100111;
   assign rom_data[6646]=8'b10000101;
   assign rom_data[6647]=8'b01100110;
   assign rom_data[6648]=8'b10000101;
   assign rom_data[6649]=8'b01100101;
   assign rom_data[6650]=8'b10000101;
   assign rom_data[6651]=8'b01100011;
   assign rom_data[6652]=8'b10000101;
   assign rom_data[6653]=8'b01100010;
   assign rom_data[6654]=8'b10000101;
   assign rom_data[6655]=8'b01100000;
   assign rom_data[6656]=8'b10000101;
   assign rom_data[6657]=8'b01011111;
   assign rom_data[6658]=8'b10000101;
   assign rom_data[6659]=8'b01011110;
   assign rom_data[6660]=8'b10000101;
   assign rom_data[6661]=8'b01011100;
   assign rom_data[6662]=8'b10000101;
   assign rom_data[6663]=8'b01011011;
   assign rom_data[6664]=8'b10000101;
   assign rom_data[6665]=8'b01011001;
   assign rom_data[6666]=8'b10000101;
   assign rom_data[6667]=8'b01011000;
   assign rom_data[6668]=8'b10000101;
   assign rom_data[6669]=8'b01010111;
   assign rom_data[6670]=8'b10000101;
   assign rom_data[6671]=8'b01010101;
   assign rom_data[6672]=8'b10000101;
   assign rom_data[6673]=8'b01010100;
   assign rom_data[6674]=8'b10000101;
   assign rom_data[6675]=8'b01010010;
   assign rom_data[6676]=8'b10000101;
   assign rom_data[6677]=8'b01010001;
   assign rom_data[6678]=8'b10000101;
   assign rom_data[6679]=8'b01010000;
   assign rom_data[6680]=8'b10000101;
   assign rom_data[6681]=8'b01001110;
   assign rom_data[6682]=8'b10000101;
   assign rom_data[6683]=8'b01001101;
   assign rom_data[6684]=8'b10000101;
   assign rom_data[6685]=8'b01001100;
   assign rom_data[6686]=8'b10000101;
   assign rom_data[6687]=8'b01001010;
   assign rom_data[6688]=8'b10000101;
   assign rom_data[6689]=8'b01001001;
   assign rom_data[6690]=8'b10000101;
   assign rom_data[6691]=8'b01001000;
   assign rom_data[6692]=8'b10000101;
   assign rom_data[6693]=8'b01000110;
   assign rom_data[6694]=8'b10000101;
   assign rom_data[6695]=8'b01000101;
   assign rom_data[6696]=8'b10000101;
   assign rom_data[6697]=8'b01000100;
   assign rom_data[6698]=8'b10000101;
   assign rom_data[6699]=8'b01000010;
   assign rom_data[6700]=8'b10000101;
   assign rom_data[6701]=8'b01000001;
   assign rom_data[6702]=8'b10000101;
   assign rom_data[6703]=8'b01000000;
   assign rom_data[6704]=8'b10000101;
   assign rom_data[6705]=8'b00111110;
   assign rom_data[6706]=8'b10000110;
   assign rom_data[6707]=8'b00111101;
   assign rom_data[6708]=8'b10000110;
   assign rom_data[6709]=8'b00111100;
   assign rom_data[6710]=8'b10000110;
   assign rom_data[6711]=8'b00111011;
   assign rom_data[6712]=8'b10000110;
   assign rom_data[6713]=8'b00111010;
   assign rom_data[6714]=8'b10000110;
   assign rom_data[6715]=8'b00111001;
   assign rom_data[6716]=8'b10000110;
   assign rom_data[6717]=8'b00111000;
   assign rom_data[6718]=8'b10000110;
   assign rom_data[6719]=8'b00110110;
   assign rom_data[6720]=8'b10000110;
   assign rom_data[6721]=8'b00110101;
   assign rom_data[6722]=8'b10000110;
   assign rom_data[6723]=8'b00110100;
   assign rom_data[6724]=8'b10000110;
   assign rom_data[6725]=8'b00110011;
   assign rom_data[6726]=8'b10000110;
   assign rom_data[6727]=8'b00110011;
   assign rom_data[6728]=8'b10000110;
   assign rom_data[6729]=8'b00110010;
   assign rom_data[6730]=8'b10000110;
   assign rom_data[6731]=8'b00110001;
   assign rom_data[6732]=8'b10000110;
   assign rom_data[6733]=8'b00110000;
   assign rom_data[6734]=8'b10000110;
   assign rom_data[6735]=8'b00101111;
   assign rom_data[6736]=8'b10000110;
   assign rom_data[6737]=8'b00101111;
   assign rom_data[6738]=8'b10000110;
   assign rom_data[6739]=8'b00101110;
   assign rom_data[6740]=8'b10000110;
   assign rom_data[6741]=8'b00101110;
   assign rom_data[6742]=8'b10000110;
   assign rom_data[6743]=8'b00101101;
   assign rom_data[6744]=8'b10000110;
   assign rom_data[6745]=8'b00101101;
   assign rom_data[6746]=8'b10000110;
   assign rom_data[6747]=8'b00101100;
   assign rom_data[6748]=8'b10000110;
   assign rom_data[6749]=8'b00101100;
   assign rom_data[6750]=8'b10000110;
   assign rom_data[6751]=8'b00101100;
   assign rom_data[6752]=8'b10000110;
   assign rom_data[6753]=8'b00101100;
   assign rom_data[6754]=8'b10000110;
   assign rom_data[6755]=8'b00101100;
   assign rom_data[6756]=8'b10000110;
   assign rom_data[6757]=8'b00101100;
   assign rom_data[6758]=8'b10000110;
   assign rom_data[6759]=8'b00101100;
   assign rom_data[6760]=8'b10000110;
   assign rom_data[6761]=8'b00101101;
   assign rom_data[6762]=8'b10000110;
   assign rom_data[6763]=8'b00101101;
   assign rom_data[6764]=8'b10000110;
   assign rom_data[6765]=8'b00101101;
   assign rom_data[6766]=8'b10000110;
   assign rom_data[6767]=8'b00101110;
   assign rom_data[6768]=8'b10000110;
   assign rom_data[6769]=8'b00101111;
   assign rom_data[6770]=8'b10000110;
   assign rom_data[6771]=8'b00101111;
   assign rom_data[6772]=8'b10000111;
   assign rom_data[6773]=8'b00110000;
   assign rom_data[6774]=8'b10000111;
   assign rom_data[6775]=8'b00110001;
   assign rom_data[6776]=8'b10000111;
   assign rom_data[6777]=8'b00110001;
   assign rom_data[6778]=8'b10000111;
   assign rom_data[6779]=8'b00110010;
   assign rom_data[6780]=8'b10000111;
   assign rom_data[6781]=8'b00110011;
   assign rom_data[6782]=8'b10000111;
   assign rom_data[6783]=8'b00110100;
   assign rom_data[6784]=8'b10000111;
   assign rom_data[6785]=8'b00110101;
   assign rom_data[6786]=8'b10000111;
   assign rom_data[6787]=8'b00110110;
   assign rom_data[6788]=8'b10000111;
   assign rom_data[6789]=8'b00110111;
   assign rom_data[6790]=8'b10000111;
   assign rom_data[6791]=8'b00111000;
   assign rom_data[6792]=8'b10000111;
   assign rom_data[6793]=8'b00111010;
   assign rom_data[6794]=8'b10000111;
   assign rom_data[6795]=8'b00111011;
   assign rom_data[6796]=8'b10000111;
   assign rom_data[6797]=8'b00111100;
   assign rom_data[6798]=8'b10000111;
   assign rom_data[6799]=8'b00111101;
   assign rom_data[6800]=8'b10000111;
   assign rom_data[6801]=8'b00111110;
   assign rom_data[6802]=8'b10000111;
   assign rom_data[6803]=8'b01000000;
   assign rom_data[6804]=8'b10000111;
   assign rom_data[6805]=8'b01000001;
   assign rom_data[6806]=8'b10000111;
   assign rom_data[6807]=8'b01000010;
   assign rom_data[6808]=8'b10000111;
   assign rom_data[6809]=8'b01000100;
   assign rom_data[6810]=8'b10000111;
   assign rom_data[6811]=8'b01000101;
   assign rom_data[6812]=8'b10000111;
   assign rom_data[6813]=8'b01000110;
   assign rom_data[6814]=8'b10000111;
   assign rom_data[6815]=8'b01001000;
   assign rom_data[6816]=8'b10000111;
   assign rom_data[6817]=8'b01001001;
   assign rom_data[6818]=8'b10000111;
   assign rom_data[6819]=8'b01001010;
   assign rom_data[6820]=8'b10000111;
   assign rom_data[6821]=8'b01001100;
   assign rom_data[6822]=8'b10000111;
   assign rom_data[6823]=8'b01001101;
   assign rom_data[6824]=8'b10000111;
   assign rom_data[6825]=8'b01001110;
   assign rom_data[6826]=8'b10000111;
   assign rom_data[6827]=8'b01010000;
   assign rom_data[6828]=8'b10000111;
   assign rom_data[6829]=8'b01010001;
   assign rom_data[6830]=8'b10000111;
   assign rom_data[6831]=8'b01010011;
   assign rom_data[6832]=8'b10000111;
   assign rom_data[6833]=8'b01010100;
   assign rom_data[6834]=8'b10000111;
   assign rom_data[6835]=8'b01010101;
   assign rom_data[6836]=8'b10000111;
   assign rom_data[6837]=8'b01010111;
   assign rom_data[6838]=8'b10000111;
   assign rom_data[6839]=8'b01011000;
   assign rom_data[6840]=8'b10000111;
   assign rom_data[6841]=8'b01011010;
   assign rom_data[6842]=8'b10000111;
   assign rom_data[6843]=8'b01011011;
   assign rom_data[6844]=8'b10000111;
   assign rom_data[6845]=8'b01011100;
   assign rom_data[6846]=8'b10000111;
   assign rom_data[6847]=8'b01011110;
   assign rom_data[6848]=8'b10000111;
   assign rom_data[6849]=8'b01011111;
   assign rom_data[6850]=8'b10000111;
   assign rom_data[6851]=8'b01100001;
   assign rom_data[6852]=8'b10001000;
   assign rom_data[6853]=8'b01100010;
   assign rom_data[6854]=8'b10001000;
   assign rom_data[6855]=8'b01100011;
   assign rom_data[6856]=8'b10001000;
   assign rom_data[6857]=8'b01100101;
   assign rom_data[6858]=8'b10001000;
   assign rom_data[6859]=8'b01100110;
   assign rom_data[6860]=8'b10001000;
   assign rom_data[6861]=8'b01101000;
   assign rom_data[6862]=8'b10001000;
   assign rom_data[6863]=8'b01101001;
   assign rom_data[6864]=8'b10001000;
   assign rom_data[6865]=8'b01101010;
   assign rom_data[6866]=8'b10001000;
   assign rom_data[6867]=8'b01101100;
   assign rom_data[6868]=8'b10001000;
   assign rom_data[6869]=8'b01101101;
   assign rom_data[6870]=8'b10001000;
   assign rom_data[6871]=8'b01101110;
   assign rom_data[6872]=8'b10001000;
   assign rom_data[6873]=8'b01110000;
   assign rom_data[6874]=8'b10001000;
   assign rom_data[6875]=8'b01110001;
   assign rom_data[6876]=8'b10001000;
   assign rom_data[6877]=8'b01110010;
   assign rom_data[6878]=8'b10001000;
   assign rom_data[6879]=8'b01110100;
   assign rom_data[6880]=8'b10001000;
   assign rom_data[6881]=8'b01110101;
   assign rom_data[6882]=8'b10001000;
   assign rom_data[6883]=8'b01110110;
   assign rom_data[6884]=8'b10001000;
   assign rom_data[6885]=8'b01110111;
   assign rom_data[6886]=8'b10001000;
   assign rom_data[6887]=8'b01111001;
   assign rom_data[6888]=8'b10001000;
   assign rom_data[6889]=8'b01111010;
   assign rom_data[6890]=8'b10001000;
   assign rom_data[6891]=8'b01111011;
   assign rom_data[6892]=8'b10001000;
   assign rom_data[6893]=8'b01111100;
   assign rom_data[6894]=8'b10001000;
   assign rom_data[6895]=8'b01111101;
   assign rom_data[6896]=8'b10001000;
   assign rom_data[6897]=8'b01111110;
   assign rom_data[6898]=8'b10001000;
   assign rom_data[6899]=8'b01111111;
   assign rom_data[6900]=8'b10001000;
   assign rom_data[6901]=8'b10000000;
   assign rom_data[6902]=8'b10001000;
   assign rom_data[6903]=8'b10000001;
   assign rom_data[6904]=8'b10001000;
   assign rom_data[6905]=8'b10000010;
   assign rom_data[6906]=8'b10001000;
   assign rom_data[6907]=8'b10000011;
   assign rom_data[6908]=8'b10001000;
   assign rom_data[6909]=8'b10000100;
   assign rom_data[6910]=8'b10001000;
   assign rom_data[6911]=8'b10000101;
   assign rom_data[6912]=8'b10001000;
   assign rom_data[6913]=8'b10000110;
   assign rom_data[6914]=8'b10001000;
   assign rom_data[6915]=8'b10000110;
   assign rom_data[6916]=8'b10001000;
   assign rom_data[6917]=8'b10000111;
   assign rom_data[6918]=8'b10001000;
   assign rom_data[6919]=8'b10001000;
   assign rom_data[6920]=8'b10001000;
   assign rom_data[6921]=8'b10001000;
   assign rom_data[6922]=8'b10001000;
   assign rom_data[6923]=8'b10001001;
   assign rom_data[6924]=8'b10001000;
   assign rom_data[6925]=8'b10001001;
   assign rom_data[6926]=8'b10001001;
   assign rom_data[6927]=8'b10001001;
   assign rom_data[6928]=8'b10001001;
   assign rom_data[6929]=8'b10001010;
   assign rom_data[6930]=8'b10001001;
   assign rom_data[6931]=8'b10001010;
   assign rom_data[6932]=8'b10001001;
   assign rom_data[6933]=8'b10001010;
   assign rom_data[6934]=8'b10001001;
   assign rom_data[6935]=8'b10001010;
   assign rom_data[6936]=8'b10001001;
   assign rom_data[6937]=8'b10001010;
   assign rom_data[6938]=8'b10001001;
   assign rom_data[6939]=8'b10001001;
   assign rom_data[6940]=8'b10001001;
   assign rom_data[6941]=8'b10001001;
   assign rom_data[6942]=8'b10001001;
   assign rom_data[6943]=8'b10001001;
   assign rom_data[6944]=8'b10001001;
   assign rom_data[6945]=8'b10001000;
   assign rom_data[6946]=8'b10001001;
   assign rom_data[6947]=8'b10001000;
   assign rom_data[6948]=8'b10001001;
   assign rom_data[6949]=8'b10000111;
   assign rom_data[6950]=8'b10001001;
   assign rom_data[6951]=8'b10000111;
   assign rom_data[6952]=8'b10001001;
   assign rom_data[6953]=8'b10000110;
   assign rom_data[6954]=8'b10001001;
   assign rom_data[6955]=8'b10000101;
   assign rom_data[6956]=8'b10001001;
   assign rom_data[6957]=8'b10000100;
   assign rom_data[6958]=8'b10001001;
   assign rom_data[6959]=8'b10000011;
   assign rom_data[6960]=8'b10001001;
   assign rom_data[6961]=8'b10000011;
   assign rom_data[6962]=8'b10001001;
   assign rom_data[6963]=8'b10000010;
   assign rom_data[6964]=8'b10001001;
   assign rom_data[6965]=8'b10000001;
   assign rom_data[6966]=8'b10001001;
   assign rom_data[6967]=8'b10000000;
   assign rom_data[6968]=8'b10001001;
   assign rom_data[6969]=8'b01111110;
   assign rom_data[6970]=8'b10001001;
   assign rom_data[6971]=8'b01111101;
   assign rom_data[6972]=8'b10001001;
   assign rom_data[6973]=8'b01111100;
   assign rom_data[6974]=8'b10001001;
   assign rom_data[6975]=8'b01111011;
   assign rom_data[6976]=8'b10001001;
   assign rom_data[6977]=8'b01111010;
   assign rom_data[6978]=8'b10001001;
   assign rom_data[6979]=8'b01111001;
   assign rom_data[6980]=8'b10001001;
   assign rom_data[6981]=8'b01110111;
   assign rom_data[6982]=8'b10001001;
   assign rom_data[6983]=8'b01110110;
   assign rom_data[6984]=8'b10001001;
   assign rom_data[6985]=8'b01110101;
   assign rom_data[6986]=8'b10001001;
   assign rom_data[6987]=8'b01110100;
   assign rom_data[6988]=8'b10001001;
   assign rom_data[6989]=8'b01110010;
   assign rom_data[6990]=8'b10001001;
   assign rom_data[6991]=8'b01110001;
   assign rom_data[6992]=8'b10001001;
   assign rom_data[6993]=8'b01110000;
   assign rom_data[6994]=8'b10001001;
   assign rom_data[6995]=8'b01101110;
   assign rom_data[6996]=8'b10001010;
   assign rom_data[6997]=8'b01101101;
   assign rom_data[6998]=8'b10001010;
   assign rom_data[6999]=8'b01101100;
   assign rom_data[7000]=8'b10001010;
   assign rom_data[7001]=8'b01101010;
   assign rom_data[7002]=8'b10001010;
   assign rom_data[7003]=8'b01101001;
   assign rom_data[7004]=8'b10001010;
   assign rom_data[7005]=8'b01100111;
   assign rom_data[7006]=8'b10001010;
   assign rom_data[7007]=8'b01100110;
   assign rom_data[7008]=8'b10001010;
   assign rom_data[7009]=8'b01100101;
   assign rom_data[7010]=8'b10001010;
   assign rom_data[7011]=8'b01100011;
   assign rom_data[7012]=8'b10001010;
   assign rom_data[7013]=8'b01100010;
   assign rom_data[7014]=8'b10001010;
   assign rom_data[7015]=8'b01100000;
   assign rom_data[7016]=8'b10001010;
   assign rom_data[7017]=8'b01011111;
   assign rom_data[7018]=8'b10001010;
   assign rom_data[7019]=8'b01011110;
   assign rom_data[7020]=8'b10001010;
   assign rom_data[7021]=8'b01011100;
   assign rom_data[7022]=8'b10001010;
   assign rom_data[7023]=8'b01011011;
   assign rom_data[7024]=8'b10001010;
   assign rom_data[7025]=8'b01011001;
   assign rom_data[7026]=8'b10001010;
   assign rom_data[7027]=8'b01011000;
   assign rom_data[7028]=8'b10001010;
   assign rom_data[7029]=8'b01010111;
   assign rom_data[7030]=8'b10001010;
   assign rom_data[7031]=8'b01010101;
   assign rom_data[7032]=8'b10001010;
   assign rom_data[7033]=8'b01010100;
   assign rom_data[7034]=8'b10001010;
   assign rom_data[7035]=8'b01010010;
   assign rom_data[7036]=8'b10001010;
   assign rom_data[7037]=8'b01010001;
   assign rom_data[7038]=8'b10001010;
   assign rom_data[7039]=8'b01010000;
   assign rom_data[7040]=8'b10001010;
   assign rom_data[7041]=8'b01001110;
   assign rom_data[7042]=8'b10001010;
   assign rom_data[7043]=8'b01001101;
   assign rom_data[7044]=8'b10001010;
   assign rom_data[7045]=8'b01001100;
   assign rom_data[7046]=8'b10001010;
   assign rom_data[7047]=8'b01001010;
   assign rom_data[7048]=8'b10001001;
   assign rom_data[7049]=8'b01001001;
   assign rom_data[7050]=8'b10001001;
   assign rom_data[7051]=8'b01001000;
   assign rom_data[7052]=8'b10001001;
   assign rom_data[7053]=8'b01000110;
   assign rom_data[7054]=8'b10001001;
   assign rom_data[7055]=8'b01000101;
   assign rom_data[7056]=8'b10001001;
   assign rom_data[7057]=8'b01000100;
   assign rom_data[7058]=8'b10001001;
   assign rom_data[7059]=8'b01000010;
   assign rom_data[7060]=8'b10001001;
   assign rom_data[7061]=8'b01000001;
   assign rom_data[7062]=8'b10001001;
   assign rom_data[7063]=8'b01000000;
   assign rom_data[7064]=8'b10001001;
   assign rom_data[7065]=8'b00111110;
   assign rom_data[7066]=8'b10001001;
   assign rom_data[7067]=8'b00111101;
   assign rom_data[7068]=8'b10001001;
   assign rom_data[7069]=8'b00111100;
   assign rom_data[7070]=8'b10001001;
   assign rom_data[7071]=8'b00111011;
   assign rom_data[7072]=8'b10001001;
   assign rom_data[7073]=8'b00111010;
   assign rom_data[7074]=8'b10001001;
   assign rom_data[7075]=8'b00111001;
   assign rom_data[7076]=8'b10001001;
   assign rom_data[7077]=8'b00111000;
   assign rom_data[7078]=8'b10001001;
   assign rom_data[7079]=8'b00110110;
   assign rom_data[7080]=8'b10001001;
   assign rom_data[7081]=8'b00110101;
   assign rom_data[7082]=8'b10001001;
   assign rom_data[7083]=8'b00110100;
   assign rom_data[7084]=8'b10001001;
   assign rom_data[7085]=8'b00110011;
   assign rom_data[7086]=8'b10001001;
   assign rom_data[7087]=8'b00110011;
   assign rom_data[7088]=8'b10001001;
   assign rom_data[7089]=8'b00110010;
   assign rom_data[7090]=8'b10001001;
   assign rom_data[7091]=8'b00110001;
   assign rom_data[7092]=8'b10001001;
   assign rom_data[7093]=8'b00110000;
   assign rom_data[7094]=8'b10001001;
   assign rom_data[7095]=8'b00101111;
   assign rom_data[7096]=8'b10001001;
   assign rom_data[7097]=8'b00101111;
   assign rom_data[7098]=8'b10001001;
   assign rom_data[7099]=8'b00101110;
   assign rom_data[7100]=8'b10001001;
   assign rom_data[7101]=8'b00101110;
   assign rom_data[7102]=8'b10001001;
   assign rom_data[7103]=8'b00101101;
   assign rom_data[7104]=8'b10001001;
   assign rom_data[7105]=8'b00101101;
   assign rom_data[7106]=8'b10001001;
   assign rom_data[7107]=8'b00101100;
   assign rom_data[7108]=8'b10001001;
   assign rom_data[7109]=8'b00101100;
   assign rom_data[7110]=8'b10001001;
   assign rom_data[7111]=8'b00101100;
   assign rom_data[7112]=8'b10001001;
   assign rom_data[7113]=8'b00101100;
   assign rom_data[7114]=8'b10001001;
   assign rom_data[7115]=8'b00101100;
   assign rom_data[7116]=8'b10001001;
   assign rom_data[7117]=8'b00101100;
   assign rom_data[7118]=8'b10001000;
   assign rom_data[7119]=8'b00101100;
   assign rom_data[7120]=8'b10001000;
   assign rom_data[7121]=8'b00101101;
   assign rom_data[7122]=8'b10001000;
   assign rom_data[7123]=8'b00101101;
   assign rom_data[7124]=8'b10001000;
   assign rom_data[7125]=8'b00101101;
   assign rom_data[7126]=8'b10001000;
   assign rom_data[7127]=8'b00101110;
   assign rom_data[7128]=8'b10001000;
   assign rom_data[7129]=8'b00101111;
   assign rom_data[7130]=8'b10001000;
   assign rom_data[7131]=8'b00101111;
   assign rom_data[7132]=8'b10001000;
   assign rom_data[7133]=8'b00110000;
   assign rom_data[7134]=8'b10001000;
   assign rom_data[7135]=8'b00110001;
   assign rom_data[7136]=8'b10001000;
   assign rom_data[7137]=8'b00110001;
   assign rom_data[7138]=8'b10001000;
   assign rom_data[7139]=8'b00110010;
   assign rom_data[7140]=8'b10001000;
   assign rom_data[7141]=8'b00110011;
   assign rom_data[7142]=8'b10001000;
   assign rom_data[7143]=8'b00110100;
   assign rom_data[7144]=8'b10001000;
   assign rom_data[7145]=8'b00110101;
   assign rom_data[7146]=8'b10001000;
   assign rom_data[7147]=8'b00110110;
   assign rom_data[7148]=8'b10001000;
   assign rom_data[7149]=8'b00110111;
   assign rom_data[7150]=8'b10001000;
   assign rom_data[7151]=8'b00111000;
   assign rom_data[7152]=8'b10001000;
   assign rom_data[7153]=8'b00111010;
   assign rom_data[7154]=8'b10001000;
   assign rom_data[7155]=8'b00111011;
   assign rom_data[7156]=8'b10001000;
   assign rom_data[7157]=8'b00111100;
   assign rom_data[7158]=8'b10001000;
   assign rom_data[7159]=8'b00111101;
   assign rom_data[7160]=8'b10001000;
   assign rom_data[7161]=8'b00111110;
   assign rom_data[7162]=8'b10001000;
   assign rom_data[7163]=8'b01000000;
   assign rom_data[7164]=8'b10001000;
   assign rom_data[7165]=8'b01000001;
   assign rom_data[7166]=8'b10001000;
   assign rom_data[7167]=8'b01000010;
   assign rom_data[7168]=8'b10001000;
   assign rom_data[7169]=8'b01000100;
   assign rom_data[7170]=8'b10001000;
   assign rom_data[7171]=8'b01000101;
   assign rom_data[7172]=8'b10001000;
   assign rom_data[7173]=8'b01000110;
   assign rom_data[7174]=8'b10001000;
   assign rom_data[7175]=8'b01001000;
   assign rom_data[7176]=8'b10001000;
   assign rom_data[7177]=8'b01001001;
   assign rom_data[7178]=8'b10001000;
   assign rom_data[7179]=8'b01001010;
   assign rom_data[7180]=8'b10001000;
   assign rom_data[7181]=8'b01001100;
   assign rom_data[7182]=8'b10001000;
   assign rom_data[7183]=8'b01001101;
   assign rom_data[7184]=8'b10001000;
   assign rom_data[7185]=8'b01001110;
   assign rom_data[7186]=8'b10001000;
   assign rom_data[7187]=8'b01010000;
   assign rom_data[7188]=8'b10001000;
   assign rom_data[7189]=8'b01010001;
   assign rom_data[7190]=8'b10001000;
   assign rom_data[7191]=8'b01010011;
   assign rom_data[7192]=8'b10000111;
   assign rom_data[7193]=8'b01010100;
   assign rom_data[7194]=8'b10000111;
   assign rom_data[7195]=8'b01010101;
   assign rom_data[7196]=8'b10000111;
   assign rom_data[7197]=8'b01010111;
   assign rom_data[7198]=8'b10000111;
   assign rom_data[7199]=8'b01011000;
   assign rom_data[7200]=8'b10000111;
   assign rom_data[7201]=8'b01011010;
   assign rom_data[7202]=8'b10000111;
   assign rom_data[7203]=8'b01011011;
   assign rom_data[7204]=8'b10000111;
   assign rom_data[7205]=8'b01011100;
   assign rom_data[7206]=8'b10000111;
   assign rom_data[7207]=8'b01011110;
   assign rom_data[7208]=8'b10000111;
   assign rom_data[7209]=8'b01011111;
   assign rom_data[7210]=8'b10000111;
   assign rom_data[7211]=8'b01100001;
   assign rom_data[7212]=8'b10000111;
   assign rom_data[7213]=8'b01100010;
   assign rom_data[7214]=8'b10000111;
   assign rom_data[7215]=8'b01100011;
   assign rom_data[7216]=8'b10000111;
   assign rom_data[7217]=8'b01100101;
   assign rom_data[7218]=8'b10000111;
   assign rom_data[7219]=8'b01100110;
   assign rom_data[7220]=8'b10000111;
   assign rom_data[7221]=8'b01101000;
   assign rom_data[7222]=8'b10000111;
   assign rom_data[7223]=8'b01101001;
   assign rom_data[7224]=8'b10000111;
   assign rom_data[7225]=8'b01101010;
   assign rom_data[7226]=8'b10000111;
   assign rom_data[7227]=8'b01101100;
   assign rom_data[7228]=8'b10000111;
   assign rom_data[7229]=8'b01101101;
   assign rom_data[7230]=8'b10000111;
   assign rom_data[7231]=8'b01101110;
   assign rom_data[7232]=8'b10000111;
   assign rom_data[7233]=8'b01110000;
   assign rom_data[7234]=8'b10000111;
   assign rom_data[7235]=8'b01110001;
   assign rom_data[7236]=8'b10000111;
   assign rom_data[7237]=8'b01110010;
   assign rom_data[7238]=8'b10000111;
   assign rom_data[7239]=8'b01110100;
   assign rom_data[7240]=8'b10000111;
   assign rom_data[7241]=8'b01110101;
   assign rom_data[7242]=8'b10000111;
   assign rom_data[7243]=8'b01110110;
   assign rom_data[7244]=8'b10000111;
   assign rom_data[7245]=8'b01110111;
   assign rom_data[7246]=8'b10000111;
   assign rom_data[7247]=8'b01111001;
   assign rom_data[7248]=8'b10000111;
   assign rom_data[7249]=8'b01111010;
   assign rom_data[7250]=8'b10000111;
   assign rom_data[7251]=8'b01111011;
   assign rom_data[7252]=8'b10000111;
   assign rom_data[7253]=8'b01111100;
   assign rom_data[7254]=8'b10000111;
   assign rom_data[7255]=8'b01111101;
   assign rom_data[7256]=8'b10000111;
   assign rom_data[7257]=8'b01111110;
   assign rom_data[7258]=8'b10000111;
   assign rom_data[7259]=8'b01111111;
   assign rom_data[7260]=8'b10000111;
   assign rom_data[7261]=8'b10000000;
   assign rom_data[7262]=8'b10000111;
   assign rom_data[7263]=8'b10000001;
   assign rom_data[7264]=8'b10000111;
   assign rom_data[7265]=8'b10000010;
   assign rom_data[7266]=8'b10000111;
   assign rom_data[7267]=8'b10000011;
   assign rom_data[7268]=8'b10000111;
   assign rom_data[7269]=8'b10000100;
   assign rom_data[7270]=8'b10000111;
   assign rom_data[7271]=8'b10000101;
   assign rom_data[7272]=8'b10000110;
   assign rom_data[7273]=8'b10000110;
   assign rom_data[7274]=8'b10000110;
   assign rom_data[7275]=8'b10000110;
   assign rom_data[7276]=8'b10000110;
   assign rom_data[7277]=8'b10000111;
   assign rom_data[7278]=8'b10000110;
   assign rom_data[7279]=8'b10001000;
   assign rom_data[7280]=8'b10000110;
   assign rom_data[7281]=8'b10001000;
   assign rom_data[7282]=8'b10000110;
   assign rom_data[7283]=8'b10001001;
   assign rom_data[7284]=8'b10000110;
   assign rom_data[7285]=8'b10001001;
   assign rom_data[7286]=8'b10000110;
   assign rom_data[7287]=8'b10001001;
   assign rom_data[7288]=8'b10000110;
   assign rom_data[7289]=8'b10001010;
   assign rom_data[7290]=8'b10000110;
   assign rom_data[7291]=8'b10001010;
   assign rom_data[7292]=8'b10000110;
   assign rom_data[7293]=8'b10001010;
   assign rom_data[7294]=8'b10000110;
   assign rom_data[7295]=8'b10001010;
   assign rom_data[7296]=8'b10000110;
   assign rom_data[7297]=8'b10001010;
   assign rom_data[7298]=8'b10000110;
   assign rom_data[7299]=8'b10001001;
   assign rom_data[7300]=8'b10000110;
   assign rom_data[7301]=8'b10001001;
   assign rom_data[7302]=8'b10000110;
   assign rom_data[7303]=8'b10001001;
   assign rom_data[7304]=8'b10000110;
   assign rom_data[7305]=8'b10001000;
   assign rom_data[7306]=8'b10000110;
   assign rom_data[7307]=8'b10001000;
   assign rom_data[7308]=8'b10000110;
   assign rom_data[7309]=8'b10000111;
   assign rom_data[7310]=8'b10000110;
   assign rom_data[7311]=8'b10000111;
   assign rom_data[7312]=8'b10000110;
   assign rom_data[7313]=8'b10000110;
   assign rom_data[7314]=8'b10000110;
   assign rom_data[7315]=8'b10000101;
   assign rom_data[7316]=8'b10000110;
   assign rom_data[7317]=8'b10000100;
   assign rom_data[7318]=8'b10000110;
   assign rom_data[7319]=8'b10000011;
   assign rom_data[7320]=8'b10000110;
   assign rom_data[7321]=8'b10000011;
   assign rom_data[7322]=8'b10000110;
   assign rom_data[7323]=8'b10000010;
   assign rom_data[7324]=8'b10000110;
   assign rom_data[7325]=8'b10000001;
   assign rom_data[7326]=8'b10000110;
   assign rom_data[7327]=8'b10000000;
   assign rom_data[7328]=8'b10000110;
   assign rom_data[7329]=8'b01111110;
   assign rom_data[7330]=8'b10000110;
   assign rom_data[7331]=8'b01111101;
   assign rom_data[7332]=8'b10000110;
   assign rom_data[7333]=8'b01111100;
   assign rom_data[7334]=8'b10000110;
   assign rom_data[7335]=8'b01111011;
   assign rom_data[7336]=8'b10000110;
   assign rom_data[7337]=8'b01111010;
   assign rom_data[7338]=8'b10000101;
   assign rom_data[7339]=8'b01111001;
   assign rom_data[7340]=8'b10000101;
   assign rom_data[7341]=8'b01110111;
   assign rom_data[7342]=8'b10000101;
   assign rom_data[7343]=8'b01110110;
   assign rom_data[7344]=8'b10000101;
   assign rom_data[7345]=8'b01110101;
   assign rom_data[7346]=8'b10000101;
   assign rom_data[7347]=8'b01110100;
   assign rom_data[7348]=8'b10000101;
   assign rom_data[7349]=8'b01110010;
   assign rom_data[7350]=8'b10000101;
   assign rom_data[7351]=8'b01110001;
   assign rom_data[7352]=8'b10000101;
   assign rom_data[7353]=8'b01110000;
   assign rom_data[7354]=8'b10000101;
   assign rom_data[7355]=8'b01101110;
   assign rom_data[7356]=8'b10000101;
   assign rom_data[7357]=8'b01101101;
   assign rom_data[7358]=8'b10000101;
   assign rom_data[7359]=8'b01101100;
   assign rom_data[7360]=8'b10000101;
   assign rom_data[7361]=8'b01101010;
   assign rom_data[7362]=8'b10000101;
   assign rom_data[7363]=8'b01101001;
   assign rom_data[7364]=8'b10000101;
   assign rom_data[7365]=8'b01100111;
   assign rom_data[7366]=8'b10000101;
   assign rom_data[7367]=8'b01100110;
   assign rom_data[7368]=8'b10000101;
   assign rom_data[7369]=8'b01100101;
   assign rom_data[7370]=8'b10000101;
   assign rom_data[7371]=8'b01100011;
   assign rom_data[7372]=8'b10000101;
   assign rom_data[7373]=8'b01100010;
   assign rom_data[7374]=8'b10000101;
   assign rom_data[7375]=8'b01100000;
   assign rom_data[7376]=8'b10000101;
   assign rom_data[7377]=8'b01011111;
   assign rom_data[7378]=8'b10000101;
   assign rom_data[7379]=8'b01011110;
   assign rom_data[7380]=8'b10000101;
   assign rom_data[7381]=8'b01011100;
   assign rom_data[7382]=8'b10000101;
   assign rom_data[7383]=8'b01011011;
   assign rom_data[7384]=8'b10000101;
   assign rom_data[7385]=8'b01011001;
   assign rom_data[7386]=8'b10000101;
   assign rom_data[7387]=8'b01011000;
   assign rom_data[7388]=8'b10000101;
   assign rom_data[7389]=8'b01010111;
   assign rom_data[7390]=8'b10000101;
   assign rom_data[7391]=8'b01010101;
   assign rom_data[7392]=8'b10000101;
   assign rom_data[7393]=8'b01010100;
   assign rom_data[7394]=8'b10000101;
   assign rom_data[7395]=8'b01010010;
   assign rom_data[7396]=8'b10000101;
   assign rom_data[7397]=8'b01010001;
   assign rom_data[7398]=8'b10000101;
   assign rom_data[7399]=8'b01010000;
   assign rom_data[7400]=8'b10000101;
   assign rom_data[7401]=8'b01001110;
   assign rom_data[7402]=8'b10000101;
   assign rom_data[7403]=8'b01001101;
   assign rom_data[7404]=8'b10000101;
   assign rom_data[7405]=8'b01001100;
   assign rom_data[7406]=8'b10000101;
   assign rom_data[7407]=8'b01001010;
   assign rom_data[7408]=8'b10000101;
   assign rom_data[7409]=8'b01001001;
   assign rom_data[7410]=8'b10000101;
   assign rom_data[7411]=8'b01001000;
   assign rom_data[7412]=8'b10000101;
   assign rom_data[7413]=8'b01000110;
   assign rom_data[7414]=8'b10000101;
   assign rom_data[7415]=8'b01000101;
   assign rom_data[7416]=8'b10000101;
   assign rom_data[7417]=8'b01000100;
   assign rom_data[7418]=8'b10000101;
   assign rom_data[7419]=8'b01000010;
   assign rom_data[7420]=8'b10000101;
   assign rom_data[7421]=8'b01000001;
   assign rom_data[7422]=8'b10000100;
   assign rom_data[7423]=8'b01000000;
   assign rom_data[7424]=8'b10000100;
   assign rom_data[7425]=8'b00111110;
   assign rom_data[7426]=8'b10000100;
   assign rom_data[7427]=8'b00111101;
   assign rom_data[7428]=8'b10000100;
   assign rom_data[7429]=8'b00111100;
   assign rom_data[7430]=8'b10000100;
   assign rom_data[7431]=8'b00111011;
   assign rom_data[7432]=8'b10000100;
   assign rom_data[7433]=8'b00111010;
   assign rom_data[7434]=8'b10000100;
   assign rom_data[7435]=8'b00111001;
   assign rom_data[7436]=8'b10000100;
   assign rom_data[7437]=8'b00111000;
   assign rom_data[7438]=8'b10000100;
   assign rom_data[7439]=8'b00110110;
   assign rom_data[7440]=8'b10000100;
   assign rom_data[7441]=8'b00110101;
   assign rom_data[7442]=8'b10000100;
   assign rom_data[7443]=8'b00110100;
   assign rom_data[7444]=8'b10000100;
   assign rom_data[7445]=8'b00110011;
   assign rom_data[7446]=8'b10000100;
   assign rom_data[7447]=8'b00110011;
   assign rom_data[7448]=8'b10000100;
   assign rom_data[7449]=8'b00110010;
   assign rom_data[7450]=8'b10000100;
   assign rom_data[7451]=8'b00110001;
   assign rom_data[7452]=8'b10000100;
   assign rom_data[7453]=8'b00110000;
   assign rom_data[7454]=8'b10000100;
   assign rom_data[7455]=8'b00101111;
   assign rom_data[7456]=8'b10000100;
   assign rom_data[7457]=8'b00101111;
   assign rom_data[7458]=8'b10000100;
   assign rom_data[7459]=8'b00101110;
   assign rom_data[7460]=8'b10000100;
   assign rom_data[7461]=8'b00101110;
   assign rom_data[7462]=8'b10000100;
   assign rom_data[7463]=8'b00101101;
   assign rom_data[7464]=8'b10000100;
   assign rom_data[7465]=8'b00101101;
   assign rom_data[7466]=8'b10000100;
   assign rom_data[7467]=8'b00101100;
   assign rom_data[7468]=8'b10000100;
   assign rom_data[7469]=8'b00101100;
   assign rom_data[7470]=8'b10000100;
   assign rom_data[7471]=8'b00101100;
   assign rom_data[7472]=8'b10000100;
   assign rom_data[7473]=8'b00101100;
   assign rom_data[7474]=8'b10000100;
   assign rom_data[7475]=8'b00101100;
   assign rom_data[7476]=8'b10000100;
   assign rom_data[7477]=8'b00101100;
   assign rom_data[7478]=8'b10000100;
   assign rom_data[7479]=8'b00101100;
   assign rom_data[7480]=8'b10000100;
   assign rom_data[7481]=8'b00101101;
   assign rom_data[7482]=8'b10000100;
   assign rom_data[7483]=8'b00101101;
   assign rom_data[7484]=8'b10000100;
   assign rom_data[7485]=8'b00101101;
   assign rom_data[7486]=8'b10000100;
   assign rom_data[7487]=8'b00101110;
   assign rom_data[7488]=8'b10000100;
   assign rom_data[7489]=8'b00101111;
   assign rom_data[7490]=8'b10000011;
   assign rom_data[7491]=8'b00101111;
   assign rom_data[7492]=8'b10000011;
   assign rom_data[7493]=8'b00110000;
   assign rom_data[7494]=8'b10000011;
   assign rom_data[7495]=8'b00110001;
   assign rom_data[7496]=8'b10000011;
   assign rom_data[7497]=8'b00110001;
   assign rom_data[7498]=8'b10000011;
   assign rom_data[7499]=8'b00110010;
   assign rom_data[7500]=8'b10000011;
   assign rom_data[7501]=8'b00110011;
   assign rom_data[7502]=8'b10000011;
   assign rom_data[7503]=8'b00110100;
   assign rom_data[7504]=8'b10000011;
   assign rom_data[7505]=8'b00110101;
   assign rom_data[7506]=8'b10000011;
   assign rom_data[7507]=8'b00110110;
   assign rom_data[7508]=8'b10000011;
   assign rom_data[7509]=8'b00110111;
   assign rom_data[7510]=8'b10000011;
   assign rom_data[7511]=8'b00111000;
   assign rom_data[7512]=8'b10000011;
   assign rom_data[7513]=8'b00111010;
   assign rom_data[7514]=8'b10000011;
   assign rom_data[7515]=8'b00111011;
   assign rom_data[7516]=8'b10000011;
   assign rom_data[7517]=8'b00111100;
   assign rom_data[7518]=8'b10000011;
   assign rom_data[7519]=8'b00111101;
   assign rom_data[7520]=8'b10000011;
   assign rom_data[7521]=8'b00111110;
   assign rom_data[7522]=8'b10000011;
   assign rom_data[7523]=8'b01000000;
   assign rom_data[7524]=8'b10000011;
   assign rom_data[7525]=8'b01000001;
   assign rom_data[7526]=8'b10000011;
   assign rom_data[7527]=8'b01000010;
   assign rom_data[7528]=8'b10000011;
   assign rom_data[7529]=8'b01000100;
   assign rom_data[7530]=8'b10000011;
   assign rom_data[7531]=8'b01000101;
   assign rom_data[7532]=8'b10000011;
   assign rom_data[7533]=8'b01000110;
   assign rom_data[7534]=8'b10000011;
   assign rom_data[7535]=8'b01001000;
   assign rom_data[7536]=8'b10000011;
   assign rom_data[7537]=8'b01001001;
   assign rom_data[7538]=8'b10000011;
   assign rom_data[7539]=8'b01001010;
   assign rom_data[7540]=8'b10000011;
   assign rom_data[7541]=8'b01001100;
   assign rom_data[7542]=8'b10000011;
   assign rom_data[7543]=8'b01001101;
   assign rom_data[7544]=8'b10000011;
   assign rom_data[7545]=8'b01001110;
   assign rom_data[7546]=8'b10000011;
   assign rom_data[7547]=8'b01010000;
   assign rom_data[7548]=8'b10000011;
   assign rom_data[7549]=8'b01010001;
   assign rom_data[7550]=8'b10000011;
   assign rom_data[7551]=8'b01010011;
   assign rom_data[7552]=8'b10000011;
   assign rom_data[7553]=8'b01010100;
   assign rom_data[7554]=8'b10000011;
   assign rom_data[7555]=8'b01010101;
   assign rom_data[7556]=8'b10000011;
   assign rom_data[7557]=8'b01010111;
   assign rom_data[7558]=8'b10000011;
   assign rom_data[7559]=8'b01011000;
   assign rom_data[7560]=8'b10000011;
   assign rom_data[7561]=8'b01011010;
   assign rom_data[7562]=8'b10000011;
   assign rom_data[7563]=8'b01011011;
   assign rom_data[7564]=8'b10000011;
   assign rom_data[7565]=8'b01011100;
   assign rom_data[7566]=8'b10000011;
   assign rom_data[7567]=8'b01011110;
   assign rom_data[7568]=8'b10000011;
   assign rom_data[7569]=8'b01011111;
   assign rom_data[7570]=8'b10000010;
   assign rom_data[7571]=8'b01100001;
   assign rom_data[7572]=8'b10000010;
   assign rom_data[7573]=8'b01100010;
   assign rom_data[7574]=8'b10000010;
   assign rom_data[7575]=8'b01100011;
   assign rom_data[7576]=8'b10000010;
   assign rom_data[7577]=8'b01100101;
   assign rom_data[7578]=8'b10000010;
   assign rom_data[7579]=8'b01100110;
   assign rom_data[7580]=8'b10000010;
   assign rom_data[7581]=8'b01101000;
   assign rom_data[7582]=8'b10000010;
   assign rom_data[7583]=8'b01101001;
   assign rom_data[7584]=8'b10000010;
   assign rom_data[7585]=8'b01101010;
   assign rom_data[7586]=8'b10000010;
   assign rom_data[7587]=8'b01101100;
   assign rom_data[7588]=8'b10000010;
   assign rom_data[7589]=8'b01101101;
   assign rom_data[7590]=8'b10000010;
   assign rom_data[7591]=8'b01101110;
   assign rom_data[7592]=8'b10000010;
   assign rom_data[7593]=8'b01110000;
   assign rom_data[7594]=8'b10000010;
   assign rom_data[7595]=8'b01110001;
   assign rom_data[7596]=8'b10000010;
   assign rom_data[7597]=8'b01110010;
   assign rom_data[7598]=8'b10000010;
   assign rom_data[7599]=8'b01110100;
   assign rom_data[7600]=8'b10000010;
   assign rom_data[7601]=8'b01110101;
   assign rom_data[7602]=8'b10000010;
   assign rom_data[7603]=8'b01110110;
   assign rom_data[7604]=8'b10000010;
   assign rom_data[7605]=8'b01110111;
   assign rom_data[7606]=8'b10000010;
   assign rom_data[7607]=8'b01111001;
   assign rom_data[7608]=8'b10000010;
   assign rom_data[7609]=8'b01111010;
   assign rom_data[7610]=8'b10000010;
   assign rom_data[7611]=8'b01111011;
   assign rom_data[7612]=8'b10000010;
   assign rom_data[7613]=8'b01111100;
   assign rom_data[7614]=8'b10000010;
   assign rom_data[7615]=8'b01111101;
   assign rom_data[7616]=8'b10000010;
   assign rom_data[7617]=8'b01111110;
   assign rom_data[7618]=8'b10000010;
   assign rom_data[7619]=8'b01111111;
   assign rom_data[7620]=8'b10000010;
   assign rom_data[7621]=8'b10000000;
   assign rom_data[7622]=8'b10000010;
   assign rom_data[7623]=8'b10000001;
   assign rom_data[7624]=8'b10000010;
   assign rom_data[7625]=8'b10000010;
   assign rom_data[7626]=8'b10000010;
   assign rom_data[7627]=8'b10000011;
   assign rom_data[7628]=8'b10000010;
   assign rom_data[7629]=8'b10000100;
   assign rom_data[7630]=8'b10000010;
   assign rom_data[7631]=8'b10000101;
   assign rom_data[7632]=8'b10000010;
   assign rom_data[7633]=8'b10000110;
   assign rom_data[7634]=8'b10000010;
   assign rom_data[7635]=8'b10000110;
   assign rom_data[7636]=8'b10000010;
   assign rom_data[7637]=8'b10000111;
   assign rom_data[7638]=8'b10000010;
   assign rom_data[7639]=8'b10001000;
   assign rom_data[7640]=8'b10000010;
   assign rom_data[7641]=8'b10001000;
   assign rom_data[7642]=8'b10000010;
   assign rom_data[7643]=8'b10001001;
   assign rom_data[7644]=8'b10000001;
   assign rom_data[7645]=8'b10001001;
   assign rom_data[7646]=8'b10000001;
   assign rom_data[7647]=8'b10001001;
   assign rom_data[7648]=8'b10000001;
   assign rom_data[7649]=8'b10001010;
   assign rom_data[7650]=8'b10000001;
   assign rom_data[7651]=8'b10001010;
   assign rom_data[7652]=8'b10000001;
   assign rom_data[7653]=8'b10001010;
   assign rom_data[7654]=8'b10000001;
   assign rom_data[7655]=8'b10001010;
   assign rom_data[7656]=8'b10000001;
   assign rom_data[7657]=8'b10001010;
   assign rom_data[7658]=8'b10000001;
   assign rom_data[7659]=8'b10001001;
   assign rom_data[7660]=8'b10000001;
   assign rom_data[7661]=8'b10001001;
   assign rom_data[7662]=8'b10000001;
   assign rom_data[7663]=8'b10001001;
   assign rom_data[7664]=8'b10000001;
   assign rom_data[7665]=8'b10001000;
   assign rom_data[7666]=8'b10000001;
   assign rom_data[7667]=8'b10001000;
   assign rom_data[7668]=8'b10000001;
   assign rom_data[7669]=8'b10000111;
   assign rom_data[7670]=8'b10000001;
   assign rom_data[7671]=8'b10000111;
   assign rom_data[7672]=8'b10000001;
   assign rom_data[7673]=8'b10000110;
   assign rom_data[7674]=8'b10000001;
   assign rom_data[7675]=8'b10000101;
   assign rom_data[7676]=8'b10000001;
   assign rom_data[7677]=8'b10000100;
   assign rom_data[7678]=8'b10000001;
   assign rom_data[7679]=8'b10000011;
   assign rom_data[7680]=8'b10000001;
   assign rom_data[7681]=8'b10000011;
   assign rom_data[7682]=8'b10000001;
   assign rom_data[7683]=8'b10000010;
   assign rom_data[7684]=8'b10000001;
   assign rom_data[7685]=8'b10000001;
   assign rom_data[7686]=8'b10000001;
   assign rom_data[7687]=8'b10000000;
   assign rom_data[7688]=8'b10000001;
   assign rom_data[7689]=8'b01111110;
   assign rom_data[7690]=8'b10000001;
   assign rom_data[7691]=8'b01111101;
   assign rom_data[7692]=8'b10000001;
   assign rom_data[7693]=8'b01111100;
   assign rom_data[7694]=8'b10000001;
   assign rom_data[7695]=8'b01111011;
   assign rom_data[7696]=8'b10000001;
   assign rom_data[7697]=8'b01111010;
   assign rom_data[7698]=8'b10000001;
   assign rom_data[7699]=8'b01111001;
   assign rom_data[7700]=8'b10000001;
   assign rom_data[7701]=8'b01110111;
   assign rom_data[7702]=8'b10000001;
   assign rom_data[7703]=8'b01110110;
   assign rom_data[7704]=8'b10000001;
   assign rom_data[7705]=8'b01110101;
   assign rom_data[7706]=8'b10000001;
   assign rom_data[7707]=8'b01110100;
   assign rom_data[7708]=8'b10000001;
   assign rom_data[7709]=8'b01110010;
   assign rom_data[7710]=8'b10000001;
   assign rom_data[7711]=8'b01110001;
   assign rom_data[7712]=8'b10000001;
   assign rom_data[7713]=8'b01110000;
   assign rom_data[7714]=8'b10000000;
   assign rom_data[7715]=8'b01101110;
   assign rom_data[7716]=8'b10000000;
   assign rom_data[7717]=8'b01101101;
   assign rom_data[7718]=8'b10000000;
   assign rom_data[7719]=8'b01101100;
   assign rom_data[7720]=8'b10000000;
   assign rom_data[7721]=8'b01101010;
   assign rom_data[7722]=8'b10000000;
   assign rom_data[7723]=8'b01101001;
   assign rom_data[7724]=8'b10000000;
   assign rom_data[7725]=8'b01100111;
   assign rom_data[7726]=8'b10000000;
   assign rom_data[7727]=8'b01100110;
   assign rom_data[7728]=8'b10000000;
   assign rom_data[7729]=8'b01100101;
   assign rom_data[7730]=8'b10000000;
   assign rom_data[7731]=8'b01100011;
   assign rom_data[7732]=8'b10000000;
   assign rom_data[7733]=8'b01100010;
   assign rom_data[7734]=8'b10000000;
   assign rom_data[7735]=8'b01100000;
   assign rom_data[7736]=8'b10000000;
   assign rom_data[7737]=8'b01011111;
   assign rom_data[7738]=8'b10000000;
   assign rom_data[7739]=8'b01011110;
   assign rom_data[7740]=8'b10000000;
   assign rom_data[7741]=8'b01011100;
   assign rom_data[7742]=8'b10000000;
   assign rom_data[7743]=8'b01011011;
   assign rom_data[7744]=8'b10000000;
   assign rom_data[7745]=8'b01011001;
   assign rom_data[7746]=8'b10000000;
   assign rom_data[7747]=8'b01011000;
   assign rom_data[7748]=8'b10000000;
   assign rom_data[7749]=8'b01010111;
   assign rom_data[7750]=8'b10000000;
   assign rom_data[7751]=8'b01010101;
   assign rom_data[7752]=8'b10000000;
   assign rom_data[7753]=8'b01010100;
   assign rom_data[7754]=8'b10000000;
   assign rom_data[7755]=8'b01010010;
   assign rom_data[7756]=8'b10000000;
   assign rom_data[7757]=8'b01010001;
   assign rom_data[7758]=8'b10000000;
   assign rom_data[7759]=8'b01010000;
   assign rom_data[7760]=8'b10000000;
   assign rom_data[7761]=8'b01001110;
   assign rom_data[7762]=8'b10000000;
   assign rom_data[7763]=8'b01001101;
   assign rom_data[7764]=8'b10000000;
   assign rom_data[7765]=8'b01001100;
   assign rom_data[7766]=8'b10000000;
   assign rom_data[7767]=8'b01001010;
   assign rom_data[7768]=8'b10000000;
   assign rom_data[7769]=8'b01001001;
   assign rom_data[7770]=8'b10000000;
   assign rom_data[7771]=8'b01001000;
   assign rom_data[7772]=8'b10000000;
   assign rom_data[7773]=8'b01000110;
   assign rom_data[7774]=8'b10000000;
   assign rom_data[7775]=8'b01000101;
   assign rom_data[7776]=8'b10000000;
   assign rom_data[7777]=8'b01000100;
   assign rom_data[7778]=8'b10000000;
   assign rom_data[7779]=8'b01000010;
   assign rom_data[7780]=8'b10000000;
   assign rom_data[7781]=8'b01000001;
   assign rom_data[7782]=8'b10000000;
   assign rom_data[7783]=8'b01000000;
   assign rom_data[7784]=8'b10000000;
   assign rom_data[7785]=8'b00111110;
   assign rom_data[7786]=8'b10000000;
   assign rom_data[7787]=8'b00111101;
   assign rom_data[7788]=8'b10000000;
   assign rom_data[7789]=8'b00111100;
   assign rom_data[7790]=8'b10000000;
   assign rom_data[7791]=8'b00111011;
   assign rom_data[7792]=8'b10000000;
   assign rom_data[7793]=8'b00111010;
   assign rom_data[7794]=8'b10000000;
   assign rom_data[7795]=8'b00111001;
   assign rom_data[7796]=8'b10000000;
   assign rom_data[7797]=8'b00111000;
   assign rom_data[7798]=8'b01111111;
   assign rom_data[7799]=8'b00110110;
   assign rom_data[7800]=8'b01111111;
   assign rom_data[7801]=8'b00110101;
   assign rom_data[7802]=8'b01111111;
   assign rom_data[7803]=8'b00110100;
   assign rom_data[7804]=8'b01111111;
   assign rom_data[7805]=8'b00110011;
   assign rom_data[7806]=8'b01111111;
   assign rom_data[7807]=8'b00110011;
   assign rom_data[7808]=8'b01111111;
   assign rom_data[7809]=8'b00110010;
   assign rom_data[7810]=8'b01111111;
   assign rom_data[7811]=8'b00110001;
   assign rom_data[7812]=8'b01111111;
   assign rom_data[7813]=8'b00110000;
   assign rom_data[7814]=8'b01111111;
   assign rom_data[7815]=8'b00101111;
   assign rom_data[7816]=8'b01111111;
   assign rom_data[7817]=8'b00101111;
   assign rom_data[7818]=8'b01111111;
   assign rom_data[7819]=8'b00101110;
   assign rom_data[7820]=8'b01111111;
   assign rom_data[7821]=8'b00101110;
   assign rom_data[7822]=8'b01111111;
   assign rom_data[7823]=8'b00101101;
   assign rom_data[7824]=8'b01111111;
   assign rom_data[7825]=8'b00101101;
   assign rom_data[7826]=8'b01111111;
   assign rom_data[7827]=8'b00101100;
   assign rom_data[7828]=8'b01111111;
   assign rom_data[7829]=8'b00101100;
   assign rom_data[7830]=8'b01111111;
   assign rom_data[7831]=8'b00101100;
   assign rom_data[7832]=8'b01111111;
   assign rom_data[7833]=8'b00101100;
   assign rom_data[7834]=8'b01111111;
   assign rom_data[7835]=8'b00101100;
   assign rom_data[7836]=8'b01111111;
   assign rom_data[7837]=8'b00101100;
   assign rom_data[7838]=8'b01111111;
   assign rom_data[7839]=8'b00101100;
   assign rom_data[7840]=8'b01111111;
   assign rom_data[7841]=8'b00101101;
   assign rom_data[7842]=8'b01111111;
   assign rom_data[7843]=8'b00101101;
   assign rom_data[7844]=8'b01111111;
   assign rom_data[7845]=8'b00101101;
   assign rom_data[7846]=8'b01111111;
   assign rom_data[7847]=8'b00101110;
   assign rom_data[7848]=8'b01111111;
   assign rom_data[7849]=8'b00101111;
   assign rom_data[7850]=8'b01111111;
   assign rom_data[7851]=8'b00101111;
   assign rom_data[7852]=8'b01111111;
   assign rom_data[7853]=8'b00110000;
   assign rom_data[7854]=8'b01111111;
   assign rom_data[7855]=8'b00110001;
   assign rom_data[7856]=8'b01111111;
   assign rom_data[7857]=8'b00110001;
   assign rom_data[7858]=8'b01111111;
   assign rom_data[7859]=8'b00110010;
   assign rom_data[7860]=8'b01111111;
   assign rom_data[7861]=8'b00110011;
   assign rom_data[7862]=8'b01111110;
   assign rom_data[7863]=8'b00110100;
   assign rom_data[7864]=8'b01111110;
   assign rom_data[7865]=8'b00110101;
   assign rom_data[7866]=8'b01111110;
   assign rom_data[7867]=8'b00110110;
   assign rom_data[7868]=8'b01111110;
   assign rom_data[7869]=8'b00110111;
   assign rom_data[7870]=8'b01111110;
   assign rom_data[7871]=8'b00111000;
   assign rom_data[7872]=8'b01111110;
   assign rom_data[7873]=8'b00111010;
   assign rom_data[7874]=8'b01111110;
   assign rom_data[7875]=8'b00111011;
   assign rom_data[7876]=8'b01111110;
   assign rom_data[7877]=8'b00111100;
   assign rom_data[7878]=8'b01111110;
   assign rom_data[7879]=8'b00111101;
   assign rom_data[7880]=8'b01111110;
   assign rom_data[7881]=8'b00111110;
   assign rom_data[7882]=8'b01111110;
   assign rom_data[7883]=8'b01000000;
   assign rom_data[7884]=8'b01111110;
   assign rom_data[7885]=8'b01000001;
   assign rom_data[7886]=8'b01111110;
   assign rom_data[7887]=8'b01000010;
   assign rom_data[7888]=8'b01111110;
   assign rom_data[7889]=8'b01000100;
   assign rom_data[7890]=8'b01111110;
   assign rom_data[7891]=8'b01000101;
   assign rom_data[7892]=8'b01111110;
   assign rom_data[7893]=8'b01000110;
   assign rom_data[7894]=8'b01111110;
   assign rom_data[7895]=8'b01001000;
   assign rom_data[7896]=8'b01111110;
   assign rom_data[7897]=8'b01001001;
   assign rom_data[7898]=8'b01111110;
   assign rom_data[7899]=8'b01001010;
   assign rom_data[7900]=8'b01111110;
   assign rom_data[7901]=8'b01001100;
   assign rom_data[7902]=8'b01111110;
   assign rom_data[7903]=8'b01001101;
   assign rom_data[7904]=8'b01111110;
   assign rom_data[7905]=8'b01001110;
   assign rom_data[7906]=8'b01111110;
   assign rom_data[7907]=8'b01010000;
   assign rom_data[7908]=8'b01111110;
   assign rom_data[7909]=8'b01010001;
   assign rom_data[7910]=8'b01111110;
   assign rom_data[7911]=8'b01010011;
   assign rom_data[7912]=8'b01111110;
   assign rom_data[7913]=8'b01010100;
   assign rom_data[7914]=8'b01111110;
   assign rom_data[7915]=8'b01010101;
   assign rom_data[7916]=8'b01111110;
   assign rom_data[7917]=8'b01010111;
   assign rom_data[7918]=8'b01111110;
   assign rom_data[7919]=8'b01011000;
   assign rom_data[7920]=8'b01111110;
   assign rom_data[7921]=8'b01011010;
   assign rom_data[7922]=8'b01111110;
   assign rom_data[7923]=8'b01011011;
   assign rom_data[7924]=8'b01111110;
   assign rom_data[7925]=8'b01011100;
   assign rom_data[7926]=8'b01111110;
   assign rom_data[7927]=8'b01011110;
   assign rom_data[7928]=8'b01111110;
   assign rom_data[7929]=8'b01011111;
   assign rom_data[7930]=8'b01111110;
   assign rom_data[7931]=8'b01100001;
   assign rom_data[7932]=8'b01111110;
   assign rom_data[7933]=8'b01100010;
   assign rom_data[7934]=8'b01111110;
   assign rom_data[7935]=8'b01100011;
   assign rom_data[7936]=8'b01111110;
   assign rom_data[7937]=8'b01100101;
   assign rom_data[7938]=8'b01111110;
   assign rom_data[7939]=8'b01100110;
   assign rom_data[7940]=8'b01111110;
   assign rom_data[7941]=8'b01101000;
   assign rom_data[7942]=8'b01111110;
   assign rom_data[7943]=8'b01101001;
   assign rom_data[7944]=8'b01111110;
   assign rom_data[7945]=8'b01101010;
   assign rom_data[7946]=8'b01111101;
   assign rom_data[7947]=8'b01101100;
   assign rom_data[7948]=8'b01111101;
   assign rom_data[7949]=8'b01101101;
   assign rom_data[7950]=8'b01111101;
   assign rom_data[7951]=8'b01101110;
   assign rom_data[7952]=8'b01111101;
   assign rom_data[7953]=8'b01110000;
   assign rom_data[7954]=8'b01111101;
   assign rom_data[7955]=8'b01110001;
   assign rom_data[7956]=8'b01111101;
   assign rom_data[7957]=8'b01110010;
   assign rom_data[7958]=8'b01111101;
   assign rom_data[7959]=8'b01110100;
   assign rom_data[7960]=8'b01111101;
   assign rom_data[7961]=8'b01110101;
   assign rom_data[7962]=8'b01111101;
   assign rom_data[7963]=8'b01110110;
   assign rom_data[7964]=8'b01111101;
   assign rom_data[7965]=8'b01110111;
   assign rom_data[7966]=8'b01111101;
   assign rom_data[7967]=8'b01111001;
   assign rom_data[7968]=8'b01111101;
   assign rom_data[7969]=8'b01111010;
   assign rom_data[7970]=8'b01111101;
   assign rom_data[7971]=8'b01111011;
   assign rom_data[7972]=8'b01111101;
   assign rom_data[7973]=8'b01111100;
   assign rom_data[7974]=8'b01111101;
   assign rom_data[7975]=8'b01111101;
   assign rom_data[7976]=8'b01111101;
   assign rom_data[7977]=8'b01111110;
   assign rom_data[7978]=8'b01111101;
   assign rom_data[7979]=8'b01111111;
   assign rom_data[7980]=8'b01111101;
   assign rom_data[7981]=8'b10000000;
   assign rom_data[7982]=8'b01111101;
   assign rom_data[7983]=8'b10000001;
   assign rom_data[7984]=8'b01111101;
   assign rom_data[7985]=8'b10000010;
   assign rom_data[7986]=8'b01111101;
   assign rom_data[7987]=8'b10000011;
   assign rom_data[7988]=8'b01111101;
   assign rom_data[7989]=8'b10000100;
   assign rom_data[7990]=8'b01111101;
   assign rom_data[7991]=8'b10000101;
   assign rom_data[7992]=8'b01111101;
   assign rom_data[7993]=8'b10000110;
   assign rom_data[7994]=8'b01111101;
   assign rom_data[7995]=8'b10000110;
   assign rom_data[7996]=8'b01111101;
   assign rom_data[7997]=8'b10000111;
   assign rom_data[7998]=8'b01111101;
   assign rom_data[7999]=8'b10001000;
   assign rom_data[8000]=8'b01111101;
   assign rom_data[8001]=8'b10001000;
   assign rom_data[8002]=8'b01111101;
   assign rom_data[8003]=8'b10001001;
   assign rom_data[8004]=8'b01111101;
   assign rom_data[8005]=8'b10001001;
   assign rom_data[8006]=8'b01111101;
   assign rom_data[8007]=8'b10001001;
   assign rom_data[8008]=8'b01111101;
   assign rom_data[8009]=8'b10001010;
   assign rom_data[8010]=8'b01111101;
   assign rom_data[8011]=8'b10001010;
   assign rom_data[8012]=8'b01111101;
   assign rom_data[8013]=8'b10001010;
   assign rom_data[8014]=8'b01111101;
   assign rom_data[8015]=8'b10001010;
   assign rom_data[8016]=8'b01111100;
   assign rom_data[8017]=8'b10001010;
   assign rom_data[8018]=8'b01111100;
   assign rom_data[8019]=8'b10001001;
   assign rom_data[8020]=8'b01111100;
   assign rom_data[8021]=8'b10001001;
   assign rom_data[8022]=8'b01111100;
   assign rom_data[8023]=8'b10001001;
   assign rom_data[8024]=8'b01111100;
   assign rom_data[8025]=8'b10001000;
   assign rom_data[8026]=8'b01111100;
   assign rom_data[8027]=8'b10001000;
   assign rom_data[8028]=8'b01111100;
   assign rom_data[8029]=8'b10000111;
   assign rom_data[8030]=8'b01111100;
   assign rom_data[8031]=8'b10000111;
   assign rom_data[8032]=8'b01111100;
   assign rom_data[8033]=8'b10000110;
   assign rom_data[8034]=8'b01111100;
   assign rom_data[8035]=8'b10000101;
   assign rom_data[8036]=8'b01111100;
   assign rom_data[8037]=8'b10000100;
   assign rom_data[8038]=8'b01111100;
   assign rom_data[8039]=8'b10000011;
   assign rom_data[8040]=8'b01111100;
   assign rom_data[8041]=8'b10000011;
   assign rom_data[8042]=8'b01111100;
   assign rom_data[8043]=8'b10000010;
   assign rom_data[8044]=8'b01111100;
   assign rom_data[8045]=8'b10000001;
   assign rom_data[8046]=8'b01111100;
   assign rom_data[8047]=8'b10000000;
   assign rom_data[8048]=8'b01111100;
   assign rom_data[8049]=8'b01111110;
   assign rom_data[8050]=8'b01111100;
   assign rom_data[8051]=8'b01111101;
   assign rom_data[8052]=8'b01111100;
   assign rom_data[8053]=8'b01111100;
   assign rom_data[8054]=8'b01111100;
   assign rom_data[8055]=8'b01111011;
   assign rom_data[8056]=8'b01111100;
   assign rom_data[8057]=8'b01111010;
   assign rom_data[8058]=8'b01111100;
   assign rom_data[8059]=8'b01111001;
   assign rom_data[8060]=8'b01111100;
   assign rom_data[8061]=8'b01110111;
   assign rom_data[8062]=8'b01111100;
   assign rom_data[8063]=8'b01110110;
   assign rom_data[8064]=8'b01111100;
   assign rom_data[8065]=8'b01110101;
   assign rom_data[8066]=8'b01111100;
   assign rom_data[8067]=8'b01110100;
   assign rom_data[8068]=8'b01111100;
   assign rom_data[8069]=8'b01110010;
   assign rom_data[8070]=8'b01111100;
   assign rom_data[8071]=8'b01110001;
   assign rom_data[8072]=8'b01111100;
   assign rom_data[8073]=8'b01110000;
   assign rom_data[8074]=8'b01111100;
   assign rom_data[8075]=8'b01101110;
   assign rom_data[8076]=8'b01111100;
   assign rom_data[8077]=8'b01101101;
   assign rom_data[8078]=8'b01111100;
   assign rom_data[8079]=8'b01101100;
   assign rom_data[8080]=8'b01111100;
   assign rom_data[8081]=8'b01101010;
   assign rom_data[8082]=8'b01111100;
   assign rom_data[8083]=8'b01101001;
   assign rom_data[8084]=8'b01111100;
   assign rom_data[8085]=8'b01100111;
   assign rom_data[8086]=8'b01111100;
   assign rom_data[8087]=8'b01100110;
   assign rom_data[8088]=8'b01111100;
   assign rom_data[8089]=8'b01100101;
   assign rom_data[8090]=8'b01111011;
   assign rom_data[8091]=8'b01100011;
   assign rom_data[8092]=8'b01111011;
   assign rom_data[8093]=8'b01100010;
   assign rom_data[8094]=8'b01111011;
   assign rom_data[8095]=8'b01100000;
   assign rom_data[8096]=8'b01111011;
   assign rom_data[8097]=8'b01011111;
   assign rom_data[8098]=8'b01111011;
   assign rom_data[8099]=8'b01011110;
   assign rom_data[8100]=8'b01111011;
   assign rom_data[8101]=8'b01011100;
   assign rom_data[8102]=8'b01111011;
   assign rom_data[8103]=8'b01011011;
   assign rom_data[8104]=8'b01111011;
   assign rom_data[8105]=8'b01011001;
   assign rom_data[8106]=8'b01111011;
   assign rom_data[8107]=8'b01011000;
   assign rom_data[8108]=8'b01111011;
   assign rom_data[8109]=8'b01010111;
   assign rom_data[8110]=8'b01111011;
   assign rom_data[8111]=8'b01010101;
   assign rom_data[8112]=8'b01111011;
   assign rom_data[8113]=8'b01010100;
   assign rom_data[8114]=8'b01111011;
   assign rom_data[8115]=8'b01010010;
   assign rom_data[8116]=8'b01111011;
   assign rom_data[8117]=8'b01010001;
   assign rom_data[8118]=8'b01111011;
   assign rom_data[8119]=8'b01010000;
   assign rom_data[8120]=8'b01111011;
   assign rom_data[8121]=8'b01001110;
   assign rom_data[8122]=8'b01111011;
   assign rom_data[8123]=8'b01001101;
   assign rom_data[8124]=8'b01111011;
   assign rom_data[8125]=8'b01001100;
   assign rom_data[8126]=8'b01111011;
   assign rom_data[8127]=8'b01001010;
   assign rom_data[8128]=8'b01111011;
   assign rom_data[8129]=8'b01001001;
   assign rom_data[8130]=8'b01111011;
   assign rom_data[8131]=8'b01001000;
   assign rom_data[8132]=8'b01111011;
   assign rom_data[8133]=8'b01000110;
   assign rom_data[8134]=8'b01111011;
   assign rom_data[8135]=8'b01000101;
   assign rom_data[8136]=8'b01111011;
   assign rom_data[8137]=8'b01000100;
   assign rom_data[8138]=8'b01111011;
   assign rom_data[8139]=8'b01000010;
   assign rom_data[8140]=8'b01111011;
   assign rom_data[8141]=8'b01000001;
   assign rom_data[8142]=8'b01111011;
   assign rom_data[8143]=8'b01000000;
   assign rom_data[8144]=8'b01111011;
   assign rom_data[8145]=8'b00111110;
   assign rom_data[8146]=8'b01111011;
   assign rom_data[8147]=8'b00111101;
   assign rom_data[8148]=8'b01111011;
   assign rom_data[8149]=8'b00111100;
   assign rom_data[8150]=8'b01111011;
   assign rom_data[8151]=8'b00111011;
   assign rom_data[8152]=8'b01111011;
   assign rom_data[8153]=8'b00111010;
   assign rom_data[8154]=8'b01111011;
   assign rom_data[8155]=8'b00111001;
   assign rom_data[8156]=8'b01111011;
   assign rom_data[8157]=8'b00111000;
   assign rom_data[8158]=8'b01111011;
   assign rom_data[8159]=8'b00110110;
   assign rom_data[8160]=8'b01111011;
   assign rom_data[8161]=8'b00110101;
   assign rom_data[8162]=8'b01111011;
   assign rom_data[8163]=8'b00110100;
   assign rom_data[8164]=8'b01111011;
   assign rom_data[8165]=8'b00110011;
   assign rom_data[8166]=8'b01111011;
   assign rom_data[8167]=8'b00110011;
   assign rom_data[8168]=8'b01111011;
   assign rom_data[8169]=8'b00110010;
   assign rom_data[8170]=8'b01111010;
   assign rom_data[8171]=8'b00110001;
   assign rom_data[8172]=8'b01111010;
   assign rom_data[8173]=8'b00110000;
   assign rom_data[8174]=8'b01111010;
   assign rom_data[8175]=8'b00101111;
   assign rom_data[8176]=8'b01111010;
   assign rom_data[8177]=8'b00101111;
   assign rom_data[8178]=8'b01111010;
   assign rom_data[8179]=8'b00101110;
   assign rom_data[8180]=8'b01111010;
   assign rom_data[8181]=8'b00101110;
   assign rom_data[8182]=8'b01111010;
   assign rom_data[8183]=8'b00101101;
   assign rom_data[8184]=8'b01111010;
   assign rom_data[8185]=8'b00101101;
   assign rom_data[8186]=8'b01111010;
   assign rom_data[8187]=8'b00101100;
   assign rom_data[8188]=8'b01111010;
   assign rom_data[8189]=8'b00101100;
   assign rom_data[8190]=8'b01111010;
   assign rom_data[8191]=8'b00101100;
   assign rom_data[8192]=8'b01111010;
   assign rom_data[8193]=8'b00101100;
   assign rom_data[8194]=8'b01111010;
   assign rom_data[8195]=8'b00101100;
   assign rom_data[8196]=8'b01111010;
   assign rom_data[8197]=8'b00101100;
   assign rom_data[8198]=8'b01111010;
   assign rom_data[8199]=8'b00101100;
   assign rom_data[8200]=8'b01111010;
   assign rom_data[8201]=8'b00101101;
   assign rom_data[8202]=8'b01111010;
   assign rom_data[8203]=8'b00101101;
   assign rom_data[8204]=8'b01111010;
   assign rom_data[8205]=8'b00101101;
   assign rom_data[8206]=8'b01111010;
   assign rom_data[8207]=8'b00101110;
   assign rom_data[8208]=8'b01111010;
   assign rom_data[8209]=8'b00101111;
   assign rom_data[8210]=8'b01111010;
   assign rom_data[8211]=8'b00101111;
   assign rom_data[8212]=8'b01111010;
   assign rom_data[8213]=8'b00110000;
   assign rom_data[8214]=8'b01111010;
   assign rom_data[8215]=8'b00110001;
   assign rom_data[8216]=8'b01111010;
   assign rom_data[8217]=8'b00110001;
   assign rom_data[8218]=8'b01111010;
   assign rom_data[8219]=8'b00110010;
   assign rom_data[8220]=8'b01111010;
   assign rom_data[8221]=8'b00110011;
   assign rom_data[8222]=8'b01111010;
   assign rom_data[8223]=8'b00110100;
   assign rom_data[8224]=8'b01111010;
   assign rom_data[8225]=8'b00110101;
   assign rom_data[8226]=8'b01111010;
   assign rom_data[8227]=8'b00110110;
   assign rom_data[8228]=8'b01111010;
   assign rom_data[8229]=8'b00110111;
   assign rom_data[8230]=8'b01111010;
   assign rom_data[8231]=8'b00111000;
   assign rom_data[8232]=8'b01111010;
   assign rom_data[8233]=8'b00111010;
   assign rom_data[8234]=8'b01111010;
   assign rom_data[8235]=8'b00111011;
   assign rom_data[8236]=8'b01111001;
   assign rom_data[8237]=8'b00111100;
   assign rom_data[8238]=8'b01111001;
   assign rom_data[8239]=8'b00111101;
   assign rom_data[8240]=8'b01111001;
   assign rom_data[8241]=8'b00111110;
   assign rom_data[8242]=8'b01111001;
   assign rom_data[8243]=8'b01000000;
   assign rom_data[8244]=8'b01111001;
   assign rom_data[8245]=8'b01000001;
   assign rom_data[8246]=8'b01111001;
   assign rom_data[8247]=8'b01000010;
   assign rom_data[8248]=8'b01111001;
   assign rom_data[8249]=8'b01000100;
   assign rom_data[8250]=8'b01111001;
   assign rom_data[8251]=8'b01000101;
   assign rom_data[8252]=8'b01111001;
   assign rom_data[8253]=8'b01000110;
   assign rom_data[8254]=8'b01111001;
   assign rom_data[8255]=8'b01001000;
   assign rom_data[8256]=8'b01111001;
   assign rom_data[8257]=8'b01001001;
   assign rom_data[8258]=8'b01111001;
   assign rom_data[8259]=8'b01001010;
   assign rom_data[8260]=8'b01111001;
   assign rom_data[8261]=8'b01001100;
   assign rom_data[8262]=8'b01111001;
   assign rom_data[8263]=8'b01001101;
   assign rom_data[8264]=8'b01111001;
   assign rom_data[8265]=8'b01001110;
   assign rom_data[8266]=8'b01111001;
   assign rom_data[8267]=8'b01010000;
   assign rom_data[8268]=8'b01111001;
   assign rom_data[8269]=8'b01010001;
   assign rom_data[8270]=8'b01111001;
   assign rom_data[8271]=8'b01010011;
   assign rom_data[8272]=8'b01111001;
   assign rom_data[8273]=8'b01010100;
   assign rom_data[8274]=8'b01111001;
   assign rom_data[8275]=8'b01010101;
   assign rom_data[8276]=8'b01111001;
   assign rom_data[8277]=8'b01010111;
   assign rom_data[8278]=8'b01111001;
   assign rom_data[8279]=8'b01011000;
   assign rom_data[8280]=8'b01111001;
   assign rom_data[8281]=8'b01011010;
   assign rom_data[8282]=8'b01111001;
   assign rom_data[8283]=8'b01011011;
   assign rom_data[8284]=8'b01111001;
   assign rom_data[8285]=8'b01011100;
   assign rom_data[8286]=8'b01111001;
   assign rom_data[8287]=8'b01011110;
   assign rom_data[8288]=8'b01111001;
   assign rom_data[8289]=8'b01011111;
   assign rom_data[8290]=8'b01111001;
   assign rom_data[8291]=8'b01100001;
   assign rom_data[8292]=8'b01111001;
   assign rom_data[8293]=8'b01100010;
   assign rom_data[8294]=8'b01111001;
   assign rom_data[8295]=8'b01100011;
   assign rom_data[8296]=8'b01111001;
   assign rom_data[8297]=8'b01100101;
   assign rom_data[8298]=8'b01111001;
   assign rom_data[8299]=8'b01100110;
   assign rom_data[8300]=8'b01111001;
   assign rom_data[8301]=8'b01101000;
   assign rom_data[8302]=8'b01111001;
   assign rom_data[8303]=8'b01101001;
   assign rom_data[8304]=8'b01111001;
   assign rom_data[8305]=8'b01101010;
   assign rom_data[8306]=8'b01111001;
   assign rom_data[8307]=8'b01101100;
   assign rom_data[8308]=8'b01111001;
   assign rom_data[8309]=8'b01101101;
   assign rom_data[8310]=8'b01111001;
   assign rom_data[8311]=8'b01101110;
   assign rom_data[8312]=8'b01111001;
   assign rom_data[8313]=8'b01110000;
   assign rom_data[8314]=8'b01111001;
   assign rom_data[8315]=8'b01110001;
   assign rom_data[8316]=8'b01111001;
   assign rom_data[8317]=8'b01110010;
   assign rom_data[8318]=8'b01111001;
   assign rom_data[8319]=8'b01110100;
   assign rom_data[8320]=8'b01111001;
   assign rom_data[8321]=8'b01110101;
   assign rom_data[8322]=8'b01111000;
   assign rom_data[8323]=8'b01110110;
   assign rom_data[8324]=8'b01111000;
   assign rom_data[8325]=8'b01110111;
   assign rom_data[8326]=8'b01111000;
   assign rom_data[8327]=8'b01111001;
   assign rom_data[8328]=8'b01111000;
   assign rom_data[8329]=8'b01111010;
   assign rom_data[8330]=8'b01111000;
   assign rom_data[8331]=8'b01111011;
   assign rom_data[8332]=8'b01111000;
   assign rom_data[8333]=8'b01111100;
   assign rom_data[8334]=8'b01111000;
   assign rom_data[8335]=8'b01111101;
   assign rom_data[8336]=8'b01111000;
   assign rom_data[8337]=8'b01111110;
   assign rom_data[8338]=8'b01111000;
   assign rom_data[8339]=8'b01111111;
   assign rom_data[8340]=8'b01111000;
   assign rom_data[8341]=8'b10000000;
   assign rom_data[8342]=8'b01111000;
   assign rom_data[8343]=8'b10000001;
   assign rom_data[8344]=8'b01111000;
   assign rom_data[8345]=8'b10000010;
   assign rom_data[8346]=8'b01111000;
   assign rom_data[8347]=8'b10000011;
   assign rom_data[8348]=8'b01111000;
   assign rom_data[8349]=8'b10000100;
   assign rom_data[8350]=8'b01111000;
   assign rom_data[8351]=8'b10000101;
   assign rom_data[8352]=8'b01111000;
   assign rom_data[8353]=8'b10000110;
   assign rom_data[8354]=8'b01111000;
   assign rom_data[8355]=8'b10000110;
   assign rom_data[8356]=8'b01111000;
   assign rom_data[8357]=8'b10000111;
   assign rom_data[8358]=8'b01111000;
   assign rom_data[8359]=8'b10001000;
   assign rom_data[8360]=8'b01111000;
   assign rom_data[8361]=8'b10001000;
   assign rom_data[8362]=8'b01111000;
   assign rom_data[8363]=8'b10001001;
   assign rom_data[8364]=8'b01111000;
   assign rom_data[8365]=8'b10001001;
   assign rom_data[8366]=8'b01111000;
   assign rom_data[8367]=8'b10001001;
   assign rom_data[8368]=8'b01111000;
   assign rom_data[8369]=8'b10001010;
   assign rom_data[8370]=8'b01111000;
   assign rom_data[8371]=8'b10001010;
   assign rom_data[8372]=8'b01111000;
   assign rom_data[8373]=8'b10001010;
   assign rom_data[8374]=8'b01111000;
   assign rom_data[8375]=8'b10001010;
   assign rom_data[8376]=8'b01111000;
   assign rom_data[8377]=8'b10001010;
   assign rom_data[8378]=8'b01111000;
   assign rom_data[8379]=8'b10001001;
   assign rom_data[8380]=8'b01111000;
   assign rom_data[8381]=8'b10001001;
   assign rom_data[8382]=8'b01111000;
   assign rom_data[8383]=8'b10001001;
   assign rom_data[8384]=8'b01111000;
   assign rom_data[8385]=8'b10001000;
   assign rom_data[8386]=8'b01111000;
   assign rom_data[8387]=8'b10001000;
   assign rom_data[8388]=8'b01110111;
   assign rom_data[8389]=8'b10000111;
   assign rom_data[8390]=8'b01110111;
   assign rom_data[8391]=8'b10000111;
   assign rom_data[8392]=8'b01110111;
   assign rom_data[8393]=8'b10000110;
   assign rom_data[8394]=8'b01110111;
   assign rom_data[8395]=8'b10000101;
   assign rom_data[8396]=8'b01110111;
   assign rom_data[8397]=8'b10000100;
   assign rom_data[8398]=8'b01110111;
   assign rom_data[8399]=8'b10000011;
   assign rom_data[8400]=8'b01110111;
   assign rom_data[8401]=8'b10000011;
   assign rom_data[8402]=8'b01110111;
   assign rom_data[8403]=8'b10000010;
   assign rom_data[8404]=8'b01110111;
   assign rom_data[8405]=8'b10000001;
   assign rom_data[8406]=8'b01110111;
   assign rom_data[8407]=8'b10000000;
   assign rom_data[8408]=8'b01110111;
   assign rom_data[8409]=8'b01111110;
   assign rom_data[8410]=8'b01110111;
   assign rom_data[8411]=8'b01111101;
   assign rom_data[8412]=8'b01110111;
   assign rom_data[8413]=8'b01111100;
   assign rom_data[8414]=8'b01110111;
   assign rom_data[8415]=8'b01111011;
   assign rom_data[8416]=8'b01110111;
   assign rom_data[8417]=8'b01111010;
   assign rom_data[8418]=8'b01110111;
   assign rom_data[8419]=8'b01111001;
   assign rom_data[8420]=8'b01110111;
   assign rom_data[8421]=8'b01110111;
   assign rom_data[8422]=8'b01110111;
   assign rom_data[8423]=8'b01110110;
   assign rom_data[8424]=8'b01110111;
   assign rom_data[8425]=8'b01110101;
   assign rom_data[8426]=8'b01110111;
   assign rom_data[8427]=8'b01110100;
   assign rom_data[8428]=8'b01110111;
   assign rom_data[8429]=8'b01110010;
   assign rom_data[8430]=8'b01110111;
   assign rom_data[8431]=8'b01110001;
   assign rom_data[8432]=8'b01110111;
   assign rom_data[8433]=8'b01110000;
   assign rom_data[8434]=8'b01110111;
   assign rom_data[8435]=8'b01101110;
   assign rom_data[8436]=8'b01110111;
   assign rom_data[8437]=8'b01101101;
   assign rom_data[8438]=8'b01110111;
   assign rom_data[8439]=8'b01101100;
   assign rom_data[8440]=8'b01110111;
   assign rom_data[8441]=8'b01101010;
   assign rom_data[8442]=8'b01110111;
   assign rom_data[8443]=8'b01101001;
   assign rom_data[8444]=8'b01110111;
   assign rom_data[8445]=8'b01100111;
   assign rom_data[8446]=8'b01110111;
   assign rom_data[8447]=8'b01100110;
   assign rom_data[8448]=8'b01110111;
   assign rom_data[8449]=8'b01100101;
   assign rom_data[8450]=8'b01110111;
   assign rom_data[8451]=8'b01100011;
   assign rom_data[8452]=8'b01110111;
   assign rom_data[8453]=8'b01100010;
   assign rom_data[8454]=8'b01110111;
   assign rom_data[8455]=8'b01100000;
   assign rom_data[8456]=8'b01110111;
   assign rom_data[8457]=8'b01011111;
   assign rom_data[8458]=8'b01110111;
   assign rom_data[8459]=8'b01011110;
   assign rom_data[8460]=8'b01110111;
   assign rom_data[8461]=8'b01011100;
   assign rom_data[8462]=8'b01110111;
   assign rom_data[8463]=8'b01011011;
   assign rom_data[8464]=8'b01110111;
   assign rom_data[8465]=8'b01011001;
   assign rom_data[8466]=8'b01110111;
   assign rom_data[8467]=8'b01011000;
   assign rom_data[8468]=8'b01110110;
   assign rom_data[8469]=8'b01010111;
   assign rom_data[8470]=8'b01110110;
   assign rom_data[8471]=8'b01010101;
   assign rom_data[8472]=8'b01110110;
   assign rom_data[8473]=8'b01010100;
   assign rom_data[8474]=8'b01110110;
   assign rom_data[8475]=8'b01010010;
   assign rom_data[8476]=8'b01110110;
   assign rom_data[8477]=8'b01010001;
   assign rom_data[8478]=8'b01110110;
   assign rom_data[8479]=8'b01010000;
   assign rom_data[8480]=8'b01110110;
   assign rom_data[8481]=8'b01001110;
   assign rom_data[8482]=8'b01110110;
   assign rom_data[8483]=8'b01001101;
   assign rom_data[8484]=8'b01110110;
   assign rom_data[8485]=8'b01001100;
   assign rom_data[8486]=8'b01110110;
   assign rom_data[8487]=8'b01001010;
   assign rom_data[8488]=8'b01110110;
   assign rom_data[8489]=8'b01001001;
   assign rom_data[8490]=8'b01110110;
   assign rom_data[8491]=8'b01001000;
   assign rom_data[8492]=8'b01110110;
   assign rom_data[8493]=8'b01000110;
   assign rom_data[8494]=8'b01110110;
   assign rom_data[8495]=8'b01000101;
   assign rom_data[8496]=8'b01110110;
   assign rom_data[8497]=8'b01000100;
   assign rom_data[8498]=8'b01110110;
   assign rom_data[8499]=8'b01000010;
   assign rom_data[8500]=8'b01110110;
   assign rom_data[8501]=8'b01000001;
   assign rom_data[8502]=8'b01110110;
   assign rom_data[8503]=8'b01000000;
   assign rom_data[8504]=8'b01110110;
   assign rom_data[8505]=8'b00111110;
   assign rom_data[8506]=8'b01110110;
   assign rom_data[8507]=8'b00111101;
   assign rom_data[8508]=8'b01110110;
   assign rom_data[8509]=8'b00111100;
   assign rom_data[8510]=8'b01110110;
   assign rom_data[8511]=8'b00111011;
   assign rom_data[8512]=8'b01110110;
   assign rom_data[8513]=8'b00111010;
   assign rom_data[8514]=8'b01110110;
   assign rom_data[8515]=8'b00111001;
   assign rom_data[8516]=8'b01110110;
   assign rom_data[8517]=8'b00111000;
   assign rom_data[8518]=8'b01110110;
   assign rom_data[8519]=8'b00110110;
   assign rom_data[8520]=8'b01110110;
   assign rom_data[8521]=8'b00110101;
   assign rom_data[8522]=8'b01110110;
   assign rom_data[8523]=8'b00110100;
   assign rom_data[8524]=8'b01110110;
   assign rom_data[8525]=8'b00110011;
   assign rom_data[8526]=8'b01110110;
   assign rom_data[8527]=8'b00110011;
   assign rom_data[8528]=8'b01110110;
   assign rom_data[8529]=8'b00110010;
   assign rom_data[8530]=8'b01110110;
   assign rom_data[8531]=8'b00110001;
   assign rom_data[8532]=8'b01110110;
   assign rom_data[8533]=8'b00110000;
   assign rom_data[8534]=8'b01110110;
   assign rom_data[8535]=8'b00101111;
   assign rom_data[8536]=8'b01110110;
   assign rom_data[8537]=8'b00101111;
   assign rom_data[8538]=8'b01110110;
   assign rom_data[8539]=8'b00101110;
   assign rom_data[8540]=8'b01110110;
   assign rom_data[8541]=8'b00101110;
   assign rom_data[8542]=8'b01110101;
   assign rom_data[8543]=8'b00101101;
   assign rom_data[8544]=8'b01110101;
   assign rom_data[8545]=8'b00101101;
   assign rom_data[8546]=8'b01110101;
   assign rom_data[8547]=8'b00101100;
   assign rom_data[8548]=8'b01110101;
   assign rom_data[8549]=8'b00101100;
   assign rom_data[8550]=8'b01110101;
   assign rom_data[8551]=8'b00101100;
   assign rom_data[8552]=8'b01110101;
   assign rom_data[8553]=8'b00101100;
   assign rom_data[8554]=8'b01110101;
   assign rom_data[8555]=8'b00101100;
   assign rom_data[8556]=8'b01110101;
   assign rom_data[8557]=8'b00101100;
   assign rom_data[8558]=8'b01110101;
   assign rom_data[8559]=8'b00101100;
   assign rom_data[8560]=8'b01110101;
   assign rom_data[8561]=8'b00101101;
   assign rom_data[8562]=8'b01110101;
   assign rom_data[8563]=8'b00101101;
   assign rom_data[8564]=8'b01110101;
   assign rom_data[8565]=8'b00101101;
   assign rom_data[8566]=8'b01110101;
   assign rom_data[8567]=8'b00101110;
   assign rom_data[8568]=8'b01110101;
   assign rom_data[8569]=8'b00101111;
   assign rom_data[8570]=8'b01110101;
   assign rom_data[8571]=8'b00101111;
   assign rom_data[8572]=8'b01110101;
   assign rom_data[8573]=8'b00110000;
   assign rom_data[8574]=8'b01110101;
   assign rom_data[8575]=8'b00110001;
   assign rom_data[8576]=8'b01110101;
   assign rom_data[8577]=8'b00110001;
   assign rom_data[8578]=8'b01110101;
   assign rom_data[8579]=8'b00110010;
   assign rom_data[8580]=8'b01110101;
   assign rom_data[8581]=8'b00110011;
   assign rom_data[8582]=8'b01110101;
   assign rom_data[8583]=8'b00110100;
   assign rom_data[8584]=8'b01110101;
   assign rom_data[8585]=8'b00110101;
   assign rom_data[8586]=8'b01110101;
   assign rom_data[8587]=8'b00110110;
   assign rom_data[8588]=8'b01110101;
   assign rom_data[8589]=8'b00110111;
   assign rom_data[8590]=8'b01110101;
   assign rom_data[8591]=8'b00111000;
   assign rom_data[8592]=8'b01110101;
   assign rom_data[8593]=8'b00111010;
   assign rom_data[8594]=8'b01110101;
   assign rom_data[8595]=8'b00111011;
   assign rom_data[8596]=8'b01110101;
   assign rom_data[8597]=8'b00111100;
   assign rom_data[8598]=8'b01110101;
   assign rom_data[8599]=8'b00111101;
   assign rom_data[8600]=8'b01110101;
   assign rom_data[8601]=8'b00111110;
   assign rom_data[8602]=8'b01110101;
   assign rom_data[8603]=8'b01000000;
   assign rom_data[8604]=8'b01110101;
   assign rom_data[8605]=8'b01000001;
   assign rom_data[8606]=8'b01110101;
   assign rom_data[8607]=8'b01000010;
   assign rom_data[8608]=8'b01110101;
   assign rom_data[8609]=8'b01000100;
   assign rom_data[8610]=8'b01110101;
   assign rom_data[8611]=8'b01000101;
   assign rom_data[8612]=8'b01110100;
   assign rom_data[8613]=8'b01000110;
   assign rom_data[8614]=8'b01110100;
   assign rom_data[8615]=8'b01001000;
   assign rom_data[8616]=8'b01110100;
   assign rom_data[8617]=8'b01001001;
   assign rom_data[8618]=8'b01110100;
   assign rom_data[8619]=8'b01001010;
   assign rom_data[8620]=8'b01110100;
   assign rom_data[8621]=8'b01001100;
   assign rom_data[8622]=8'b01110100;
   assign rom_data[8623]=8'b01001101;
   assign rom_data[8624]=8'b01110100;
   assign rom_data[8625]=8'b01001110;
   assign rom_data[8626]=8'b01110100;
   assign rom_data[8627]=8'b01010000;
   assign rom_data[8628]=8'b01110100;
   assign rom_data[8629]=8'b01010001;
   assign rom_data[8630]=8'b01110100;
   assign rom_data[8631]=8'b01010011;
   assign rom_data[8632]=8'b01110100;
   assign rom_data[8633]=8'b01010100;
   assign rom_data[8634]=8'b01110100;
   assign rom_data[8635]=8'b01010101;
   assign rom_data[8636]=8'b01110100;
   assign rom_data[8637]=8'b01010111;
   assign rom_data[8638]=8'b01110100;
   assign rom_data[8639]=8'b01011000;
   assign rom_data[8640]=8'b01110100;
   assign rom_data[8641]=8'b01011010;
   assign rom_data[8642]=8'b01110100;
   assign rom_data[8643]=8'b01011011;
   assign rom_data[8644]=8'b01110100;
   assign rom_data[8645]=8'b01011100;
   assign rom_data[8646]=8'b01110100;
   assign rom_data[8647]=8'b01011110;
   assign rom_data[8648]=8'b01110100;
   assign rom_data[8649]=8'b01011111;
   assign rom_data[8650]=8'b01110100;
   assign rom_data[8651]=8'b01100001;
   assign rom_data[8652]=8'b01110100;
   assign rom_data[8653]=8'b01100010;
   assign rom_data[8654]=8'b01110100;
   assign rom_data[8655]=8'b01100011;
   assign rom_data[8656]=8'b01110100;
   assign rom_data[8657]=8'b01100101;
   assign rom_data[8658]=8'b01110100;
   assign rom_data[8659]=8'b01100110;
   assign rom_data[8660]=8'b01110100;
   assign rom_data[8661]=8'b01101000;
   assign rom_data[8662]=8'b01110100;
   assign rom_data[8663]=8'b01101001;
   assign rom_data[8664]=8'b01110100;
   assign rom_data[8665]=8'b01101010;
   assign rom_data[8666]=8'b01110100;
   assign rom_data[8667]=8'b01101100;
   assign rom_data[8668]=8'b01110100;
   assign rom_data[8669]=8'b01101101;
   assign rom_data[8670]=8'b01110100;
   assign rom_data[8671]=8'b01101110;
   assign rom_data[8672]=8'b01110100;
   assign rom_data[8673]=8'b01110000;
   assign rom_data[8674]=8'b01110100;
   assign rom_data[8675]=8'b01110001;
   assign rom_data[8676]=8'b01110100;
   assign rom_data[8677]=8'b01110010;
   assign rom_data[8678]=8'b01110100;
   assign rom_data[8679]=8'b01110100;
   assign rom_data[8680]=8'b01110100;
   assign rom_data[8681]=8'b01110101;
   assign rom_data[8682]=8'b01110100;
   assign rom_data[8683]=8'b01110110;
   assign rom_data[8684]=8'b01110100;
   assign rom_data[8685]=8'b01110111;
   assign rom_data[8686]=8'b01110100;
   assign rom_data[8687]=8'b01111001;
   assign rom_data[8688]=8'b01110100;
   assign rom_data[8689]=8'b01111010;
   assign rom_data[8690]=8'b01110100;
   assign rom_data[8691]=8'b01111011;
   assign rom_data[8692]=8'b01110100;
   assign rom_data[8693]=8'b01111100;
   assign rom_data[8694]=8'b01110100;
   assign rom_data[8695]=8'b01111101;
   assign rom_data[8696]=8'b01110011;
   assign rom_data[8697]=8'b01111110;
   assign rom_data[8698]=8'b01110011;
   assign rom_data[8699]=8'b01111111;
   assign rom_data[8700]=8'b01110011;
   assign rom_data[8701]=8'b10000000;
   assign rom_data[8702]=8'b01110011;
   assign rom_data[8703]=8'b10000001;
   assign rom_data[8704]=8'b01110011;
   assign rom_data[8705]=8'b10000010;
   assign rom_data[8706]=8'b01110011;
   assign rom_data[8707]=8'b10000011;
   assign rom_data[8708]=8'b01110011;
   assign rom_data[8709]=8'b10000100;
   assign rom_data[8710]=8'b01110011;
   assign rom_data[8711]=8'b10000101;
   assign rom_data[8712]=8'b01110011;
   assign rom_data[8713]=8'b10000110;
   assign rom_data[8714]=8'b01110011;
   assign rom_data[8715]=8'b10000110;
   assign rom_data[8716]=8'b01110011;
   assign rom_data[8717]=8'b10000111;
   assign rom_data[8718]=8'b01110011;
   assign rom_data[8719]=8'b10001000;
   assign rom_data[8720]=8'b01110011;
   assign rom_data[8721]=8'b10001000;
   assign rom_data[8722]=8'b01110011;
   assign rom_data[8723]=8'b10001001;
   assign rom_data[8724]=8'b01110011;
   assign rom_data[8725]=8'b10001001;
   assign rom_data[8726]=8'b01110011;
   assign rom_data[8727]=8'b10001001;
   assign rom_data[8728]=8'b01110011;
   assign rom_data[8729]=8'b10001010;
   assign rom_data[8730]=8'b01110011;
   assign rom_data[8731]=8'b10001010;
   assign rom_data[8732]=8'b01110011;
   assign rom_data[8733]=8'b10001010;
   assign rom_data[8734]=8'b01110011;
   assign rom_data[8735]=8'b10001010;
   assign rom_data[8736]=8'b01110011;
   assign rom_data[8737]=8'b10001010;
   assign rom_data[8738]=8'b01110011;
   assign rom_data[8739]=8'b10001001;
   assign rom_data[8740]=8'b01110011;
   assign rom_data[8741]=8'b10001001;
   assign rom_data[8742]=8'b01110011;
   assign rom_data[8743]=8'b10001001;
   assign rom_data[8744]=8'b01110011;
   assign rom_data[8745]=8'b10001000;
   assign rom_data[8746]=8'b01110011;
   assign rom_data[8747]=8'b10001000;
   assign rom_data[8748]=8'b01110011;
   assign rom_data[8749]=8'b10000111;
   assign rom_data[8750]=8'b01110011;
   assign rom_data[8751]=8'b10000111;
   assign rom_data[8752]=8'b01110011;
   assign rom_data[8753]=8'b10000110;
   assign rom_data[8754]=8'b01110011;
   assign rom_data[8755]=8'b10000101;
   assign rom_data[8756]=8'b01110011;
   assign rom_data[8757]=8'b10000100;
   assign rom_data[8758]=8'b01110011;
   assign rom_data[8759]=8'b10000011;
   assign rom_data[8760]=8'b01110010;
   assign rom_data[8761]=8'b10000011;
   assign rom_data[8762]=8'b01110010;
   assign rom_data[8763]=8'b10000010;
   assign rom_data[8764]=8'b01110010;
   assign rom_data[8765]=8'b10000001;
   assign rom_data[8766]=8'b01110010;
   assign rom_data[8767]=8'b10000000;
   assign rom_data[8768]=8'b01110010;
   assign rom_data[8769]=8'b01111110;
   assign rom_data[8770]=8'b01110010;
   assign rom_data[8771]=8'b01111101;
   assign rom_data[8772]=8'b01110010;
   assign rom_data[8773]=8'b01111100;
   assign rom_data[8774]=8'b01110010;
   assign rom_data[8775]=8'b01111011;
   assign rom_data[8776]=8'b01110010;
   assign rom_data[8777]=8'b01111010;
   assign rom_data[8778]=8'b01110010;
   assign rom_data[8779]=8'b01111001;
   assign rom_data[8780]=8'b01110010;
   assign rom_data[8781]=8'b01110111;
   assign rom_data[8782]=8'b01110010;
   assign rom_data[8783]=8'b01110110;
   assign rom_data[8784]=8'b01110010;
   assign rom_data[8785]=8'b01110101;
   assign rom_data[8786]=8'b01110010;
   assign rom_data[8787]=8'b01110100;
   assign rom_data[8788]=8'b01110010;
   assign rom_data[8789]=8'b01110010;
   assign rom_data[8790]=8'b01110010;
   assign rom_data[8791]=8'b01110001;
   assign rom_data[8792]=8'b01110010;
   assign rom_data[8793]=8'b01110000;
   assign rom_data[8794]=8'b01110010;
   assign rom_data[8795]=8'b01101110;
   assign rom_data[8796]=8'b01110010;
   assign rom_data[8797]=8'b01101101;
   assign rom_data[8798]=8'b01110010;
   assign rom_data[8799]=8'b01101100;
   assign rom_data[8800]=8'b01110010;
   assign rom_data[8801]=8'b01101010;
   assign rom_data[8802]=8'b01110010;
   assign rom_data[8803]=8'b01101001;
   assign rom_data[8804]=8'b01110010;
   assign rom_data[8805]=8'b01100111;
   assign rom_data[8806]=8'b01110010;
   assign rom_data[8807]=8'b01100110;
   assign rom_data[8808]=8'b01110010;
   assign rom_data[8809]=8'b01100101;
   assign rom_data[8810]=8'b01110010;
   assign rom_data[8811]=8'b01100011;
   assign rom_data[8812]=8'b01110010;
   assign rom_data[8813]=8'b01100010;
   assign rom_data[8814]=8'b01110010;
   assign rom_data[8815]=8'b01100000;
   assign rom_data[8816]=8'b01110010;
   assign rom_data[8817]=8'b01011111;
   assign rom_data[8818]=8'b01110010;
   assign rom_data[8819]=8'b01011110;
   assign rom_data[8820]=8'b01110010;
   assign rom_data[8821]=8'b01011100;
   assign rom_data[8822]=8'b01110010;
   assign rom_data[8823]=8'b01011011;
   assign rom_data[8824]=8'b01110010;
   assign rom_data[8825]=8'b01011001;
   assign rom_data[8826]=8'b01110010;
   assign rom_data[8827]=8'b01011000;
   assign rom_data[8828]=8'b01110010;
   assign rom_data[8829]=8'b01010111;
   assign rom_data[8830]=8'b01110010;
   assign rom_data[8831]=8'b01010101;
   assign rom_data[8832]=8'b01110010;
   assign rom_data[8833]=8'b01010100;
   assign rom_data[8834]=8'b01110010;
   assign rom_data[8835]=8'b01010010;
   assign rom_data[8836]=8'b01110010;
   assign rom_data[8837]=8'b01010001;
   assign rom_data[8838]=8'b01110010;
   assign rom_data[8839]=8'b01010000;
   assign rom_data[8840]=8'b01110010;
   assign rom_data[8841]=8'b01001110;
   assign rom_data[8842]=8'b01110010;
   assign rom_data[8843]=8'b01001101;
   assign rom_data[8844]=8'b01110001;
   assign rom_data[8845]=8'b01001100;
   assign rom_data[8846]=8'b01110001;
   assign rom_data[8847]=8'b01001010;
   assign rom_data[8848]=8'b01110001;
   assign rom_data[8849]=8'b01001001;
   assign rom_data[8850]=8'b01110001;
   assign rom_data[8851]=8'b01001000;
   assign rom_data[8852]=8'b01110001;
   assign rom_data[8853]=8'b01000110;
   assign rom_data[8854]=8'b01110001;
   assign rom_data[8855]=8'b01000101;
   assign rom_data[8856]=8'b01110001;
   assign rom_data[8857]=8'b01000100;
   assign rom_data[8858]=8'b01110001;
   assign rom_data[8859]=8'b01000010;
   assign rom_data[8860]=8'b01110001;
   assign rom_data[8861]=8'b01000001;
   assign rom_data[8862]=8'b01110001;
   assign rom_data[8863]=8'b01000000;
   assign rom_data[8864]=8'b01110001;
   assign rom_data[8865]=8'b00111110;
   assign rom_data[8866]=8'b01110001;
   assign rom_data[8867]=8'b00111101;
   assign rom_data[8868]=8'b01110001;
   assign rom_data[8869]=8'b00111100;
   assign rom_data[8870]=8'b01110001;
   assign rom_data[8871]=8'b00111011;
   assign rom_data[8872]=8'b01110001;
   assign rom_data[8873]=8'b00111010;
   assign rom_data[8874]=8'b01110001;
   assign rom_data[8875]=8'b00111001;
   assign rom_data[8876]=8'b01110001;
   assign rom_data[8877]=8'b00110111;
   assign rom_data[8878]=8'b01110001;
   assign rom_data[8879]=8'b00110110;
   assign rom_data[8880]=8'b01110001;
   assign rom_data[8881]=8'b00110101;
   assign rom_data[8882]=8'b01110001;
   assign rom_data[8883]=8'b00110100;
   assign rom_data[8884]=8'b01110001;
   assign rom_data[8885]=8'b00110011;
   assign rom_data[8886]=8'b01110001;
   assign rom_data[8887]=8'b00110011;
   assign rom_data[8888]=8'b01110001;
   assign rom_data[8889]=8'b00110010;
   assign rom_data[8890]=8'b01110001;
   assign rom_data[8891]=8'b00110001;
   assign rom_data[8892]=8'b01110001;
   assign rom_data[8893]=8'b00110000;
   assign rom_data[8894]=8'b01110001;
   assign rom_data[8895]=8'b00101111;
   assign rom_data[8896]=8'b01110001;
   assign rom_data[8897]=8'b00101111;
   assign rom_data[8898]=8'b01110001;
   assign rom_data[8899]=8'b00101110;
   assign rom_data[8900]=8'b01110001;
   assign rom_data[8901]=8'b00101110;
   assign rom_data[8902]=8'b01110001;
   assign rom_data[8903]=8'b00101101;
   assign rom_data[8904]=8'b01110001;
   assign rom_data[8905]=8'b00101101;
   assign rom_data[8906]=8'b01110001;
   assign rom_data[8907]=8'b00101100;
   assign rom_data[8908]=8'b01110001;
   assign rom_data[8909]=8'b00101100;
   assign rom_data[8910]=8'b01110001;
   assign rom_data[8911]=8'b00101100;
   assign rom_data[8912]=8'b01110001;
   assign rom_data[8913]=8'b00101100;
   assign rom_data[8914]=8'b01110000;
   assign rom_data[8915]=8'b00101100;
   assign rom_data[8916]=8'b01110000;
   assign rom_data[8917]=8'b00101100;
   assign rom_data[8918]=8'b01110000;
   assign rom_data[8919]=8'b00101100;
   assign rom_data[8920]=8'b01110000;
   assign rom_data[8921]=8'b00101101;
   assign rom_data[8922]=8'b01110000;
   assign rom_data[8923]=8'b00101101;
   assign rom_data[8924]=8'b01110000;
   assign rom_data[8925]=8'b00101101;
   assign rom_data[8926]=8'b01110000;
   assign rom_data[8927]=8'b00101110;
   assign rom_data[8928]=8'b01110000;
   assign rom_data[8929]=8'b00101111;
   assign rom_data[8930]=8'b01110000;
   assign rom_data[8931]=8'b00101111;
   assign rom_data[8932]=8'b01110000;
   assign rom_data[8933]=8'b00110000;
   assign rom_data[8934]=8'b01110000;
   assign rom_data[8935]=8'b00110001;
   assign rom_data[8936]=8'b01110000;
   assign rom_data[8937]=8'b00110001;
   assign rom_data[8938]=8'b01110000;
   assign rom_data[8939]=8'b00110010;
   assign rom_data[8940]=8'b01110000;
   assign rom_data[8941]=8'b00110011;
   assign rom_data[8942]=8'b01110000;
   assign rom_data[8943]=8'b00110100;
   assign rom_data[8944]=8'b01110000;
   assign rom_data[8945]=8'b00110101;
   assign rom_data[8946]=8'b01110000;
   assign rom_data[8947]=8'b00110110;
   assign rom_data[8948]=8'b01110000;
   assign rom_data[8949]=8'b00110111;
   assign rom_data[8950]=8'b01110000;
   assign rom_data[8951]=8'b00111000;
   assign rom_data[8952]=8'b01110000;
   assign rom_data[8953]=8'b00111010;
   assign rom_data[8954]=8'b01110000;
   assign rom_data[8955]=8'b00111011;
   assign rom_data[8956]=8'b01110000;
   assign rom_data[8957]=8'b00111100;
   assign rom_data[8958]=8'b01110000;
   assign rom_data[8959]=8'b00111101;
   assign rom_data[8960]=8'b01110000;
   assign rom_data[8961]=8'b00111110;
   assign rom_data[8962]=8'b01110000;
   assign rom_data[8963]=8'b01000000;
   assign rom_data[8964]=8'b01110000;
   assign rom_data[8965]=8'b01000001;
   assign rom_data[8966]=8'b01110000;
   assign rom_data[8967]=8'b01000010;
   assign rom_data[8968]=8'b01110000;
   assign rom_data[8969]=8'b01000100;
   assign rom_data[8970]=8'b01110000;
   assign rom_data[8971]=8'b01000101;
   assign rom_data[8972]=8'b01110000;
   assign rom_data[8973]=8'b01000110;
   assign rom_data[8974]=8'b01110000;
   assign rom_data[8975]=8'b01001000;
   assign rom_data[8976]=8'b01110000;
   assign rom_data[8977]=8'b01001001;
   assign rom_data[8978]=8'b01110000;
   assign rom_data[8979]=8'b01001010;
   assign rom_data[8980]=8'b01110000;
   assign rom_data[8981]=8'b01001100;
   assign rom_data[8982]=8'b01110000;
   assign rom_data[8983]=8'b01001101;
   assign rom_data[8984]=8'b01110000;
   assign rom_data[8985]=8'b01001110;
   assign rom_data[8986]=8'b01110000;
   assign rom_data[8987]=8'b01010000;
   assign rom_data[8988]=8'b01101111;
   assign rom_data[8989]=8'b01010001;
   assign rom_data[8990]=8'b01101111;
   assign rom_data[8991]=8'b01010011;
   assign rom_data[8992]=8'b01101111;
   assign rom_data[8993]=8'b01010100;
   assign rom_data[8994]=8'b01101111;
   assign rom_data[8995]=8'b01010101;
   assign rom_data[8996]=8'b01101111;
   assign rom_data[8997]=8'b01010111;
   assign rom_data[8998]=8'b01101111;
   assign rom_data[8999]=8'b01011000;
   assign rom_data[9000]=8'b01101111;
   assign rom_data[9001]=8'b01011010;
   assign rom_data[9002]=8'b01101111;
   assign rom_data[9003]=8'b01011011;
   assign rom_data[9004]=8'b01101111;
   assign rom_data[9005]=8'b01011100;
   assign rom_data[9006]=8'b01101111;
   assign rom_data[9007]=8'b01011110;
   assign rom_data[9008]=8'b01101111;
   assign rom_data[9009]=8'b01011111;
   assign rom_data[9010]=8'b01101111;
   assign rom_data[9011]=8'b01100001;
   assign rom_data[9012]=8'b01101111;
   assign rom_data[9013]=8'b01100010;
   assign rom_data[9014]=8'b01101111;
   assign rom_data[9015]=8'b01100011;
   assign rom_data[9016]=8'b01101111;
   assign rom_data[9017]=8'b01100101;
   assign rom_data[9018]=8'b01101111;
   assign rom_data[9019]=8'b01100110;
   assign rom_data[9020]=8'b01101111;
   assign rom_data[9021]=8'b01101000;
   assign rom_data[9022]=8'b01101111;
   assign rom_data[9023]=8'b01101001;
   assign rom_data[9024]=8'b01101111;
   assign rom_data[9025]=8'b01101010;
   assign rom_data[9026]=8'b01101111;
   assign rom_data[9027]=8'b01101100;
   assign rom_data[9028]=8'b01101111;
   assign rom_data[9029]=8'b01101101;
   assign rom_data[9030]=8'b01101111;
   assign rom_data[9031]=8'b01101110;
   assign rom_data[9032]=8'b01101111;
   assign rom_data[9033]=8'b01110000;
   assign rom_data[9034]=8'b01101111;
   assign rom_data[9035]=8'b01110001;
   assign rom_data[9036]=8'b01101111;
   assign rom_data[9037]=8'b01110010;
   assign rom_data[9038]=8'b01101111;
   assign rom_data[9039]=8'b01110100;
   assign rom_data[9040]=8'b01101111;
   assign rom_data[9041]=8'b01110101;
   assign rom_data[9042]=8'b01101111;
   assign rom_data[9043]=8'b01110110;
   assign rom_data[9044]=8'b01101111;
   assign rom_data[9045]=8'b01110111;
   assign rom_data[9046]=8'b01101111;
   assign rom_data[9047]=8'b01111001;
   assign rom_data[9048]=8'b01101111;
   assign rom_data[9049]=8'b01111010;
   assign rom_data[9050]=8'b01101111;
   assign rom_data[9051]=8'b01111011;
   assign rom_data[9052]=8'b01101111;
   assign rom_data[9053]=8'b01111100;
   assign rom_data[9054]=8'b01101111;
   assign rom_data[9055]=8'b01111101;
   assign rom_data[9056]=8'b01101111;
   assign rom_data[9057]=8'b01111110;
   assign rom_data[9058]=8'b01101111;
   assign rom_data[9059]=8'b01111111;
   assign rom_data[9060]=8'b01101111;
   assign rom_data[9061]=8'b10000000;
   assign rom_data[9062]=8'b01101111;
   assign rom_data[9063]=8'b10000001;
   assign rom_data[9064]=8'b01101111;
   assign rom_data[9065]=8'b10000010;
   assign rom_data[9066]=8'b01101111;
   assign rom_data[9067]=8'b10000011;
   assign rom_data[9068]=8'b01101110;
   assign rom_data[9069]=8'b10000100;
   assign rom_data[9070]=8'b01101110;
   assign rom_data[9071]=8'b10000101;
   assign rom_data[9072]=8'b01101110;
   assign rom_data[9073]=8'b10000110;
   assign rom_data[9074]=8'b01101110;
   assign rom_data[9075]=8'b10000110;
   assign rom_data[9076]=8'b01101110;
   assign rom_data[9077]=8'b10000111;
   assign rom_data[9078]=8'b01101110;
   assign rom_data[9079]=8'b10001000;
   assign rom_data[9080]=8'b01101110;
   assign rom_data[9081]=8'b10001000;
   assign rom_data[9082]=8'b01101110;
   assign rom_data[9083]=8'b10001001;
   assign rom_data[9084]=8'b01101110;
   assign rom_data[9085]=8'b10001001;
   assign rom_data[9086]=8'b01101110;
   assign rom_data[9087]=8'b10001001;
   assign rom_data[9088]=8'b01101110;
   assign rom_data[9089]=8'b10001010;
   assign rom_data[9090]=8'b01101110;
   assign rom_data[9091]=8'b10001010;
   assign rom_data[9092]=8'b01101110;
   assign rom_data[9093]=8'b10001010;
   assign rom_data[9094]=8'b01101110;
   assign rom_data[9095]=8'b10001010;
   assign rom_data[9096]=8'b01101110;
   assign rom_data[9097]=8'b10001010;
   assign rom_data[9098]=8'b01101110;
   assign rom_data[9099]=8'b10001001;
   assign rom_data[9100]=8'b01101110;
   assign rom_data[9101]=8'b10001001;
   assign rom_data[9102]=8'b01101110;
   assign rom_data[9103]=8'b10001001;
   assign rom_data[9104]=8'b01101110;
   assign rom_data[9105]=8'b10001000;
   assign rom_data[9106]=8'b01101110;
   assign rom_data[9107]=8'b10001000;
   assign rom_data[9108]=8'b01101110;
   assign rom_data[9109]=8'b10000111;
   assign rom_data[9110]=8'b01101110;
   assign rom_data[9111]=8'b10000111;
   assign rom_data[9112]=8'b01101110;
   assign rom_data[9113]=8'b10000110;
   assign rom_data[9114]=8'b01101110;
   assign rom_data[9115]=8'b10000101;
   assign rom_data[9116]=8'b01101110;
   assign rom_data[9117]=8'b10000100;
   assign rom_data[9118]=8'b01101110;
   assign rom_data[9119]=8'b10000011;
   assign rom_data[9120]=8'b01101110;
   assign rom_data[9121]=8'b10000011;
   assign rom_data[9122]=8'b01101110;
   assign rom_data[9123]=8'b10000010;
   assign rom_data[9124]=8'b01101110;
   assign rom_data[9125]=8'b10000001;
   assign rom_data[9126]=8'b01101110;
   assign rom_data[9127]=8'b10000000;
   assign rom_data[9128]=8'b01101110;
   assign rom_data[9129]=8'b01111110;
   assign rom_data[9130]=8'b01101110;
   assign rom_data[9131]=8'b01111101;
   assign rom_data[9132]=8'b01101110;
   assign rom_data[9133]=8'b01111100;
   assign rom_data[9134]=8'b01101110;
   assign rom_data[9135]=8'b01111011;
   assign rom_data[9136]=8'b01101101;
   assign rom_data[9137]=8'b01111010;
   assign rom_data[9138]=8'b01101101;
   assign rom_data[9139]=8'b01111001;
   assign rom_data[9140]=8'b01101101;
   assign rom_data[9141]=8'b01110111;
   assign rom_data[9142]=8'b01101101;
   assign rom_data[9143]=8'b01110110;
   assign rom_data[9144]=8'b01101101;
   assign rom_data[9145]=8'b01110101;
   assign rom_data[9146]=8'b01101101;
   assign rom_data[9147]=8'b01110100;
   assign rom_data[9148]=8'b01101101;
   assign rom_data[9149]=8'b01110010;
   assign rom_data[9150]=8'b01101101;
   assign rom_data[9151]=8'b01110001;
   assign rom_data[9152]=8'b01101101;
   assign rom_data[9153]=8'b01110000;
   assign rom_data[9154]=8'b01101101;
   assign rom_data[9155]=8'b01101110;
   assign rom_data[9156]=8'b01101101;
   assign rom_data[9157]=8'b01101101;
   assign rom_data[9158]=8'b01101101;
   assign rom_data[9159]=8'b01101100;
   assign rom_data[9160]=8'b01101101;
   assign rom_data[9161]=8'b01101010;
   assign rom_data[9162]=8'b01101101;
   assign rom_data[9163]=8'b01101001;
   assign rom_data[9164]=8'b01101101;
   assign rom_data[9165]=8'b01100111;
   assign rom_data[9166]=8'b01101101;
   assign rom_data[9167]=8'b01100110;
   assign rom_data[9168]=8'b01101101;
   assign rom_data[9169]=8'b01100101;
   assign rom_data[9170]=8'b01101101;
   assign rom_data[9171]=8'b01100011;
   assign rom_data[9172]=8'b01101101;
   assign rom_data[9173]=8'b01100010;
   assign rom_data[9174]=8'b01101101;
   assign rom_data[9175]=8'b01100000;
   assign rom_data[9176]=8'b01101101;
   assign rom_data[9177]=8'b01011111;
   assign rom_data[9178]=8'b01101101;
   assign rom_data[9179]=8'b01011110;
   assign rom_data[9180]=8'b01101101;
   assign rom_data[9181]=8'b01011100;
   assign rom_data[9182]=8'b01101101;
   assign rom_data[9183]=8'b01011011;
   assign rom_data[9184]=8'b01101101;
   assign rom_data[9185]=8'b01011001;
   assign rom_data[9186]=8'b01101101;
   assign rom_data[9187]=8'b01011000;
   assign rom_data[9188]=8'b01101101;
   assign rom_data[9189]=8'b01010111;
   assign rom_data[9190]=8'b01101101;
   assign rom_data[9191]=8'b01010101;
   assign rom_data[9192]=8'b01101101;
   assign rom_data[9193]=8'b01010100;
   assign rom_data[9194]=8'b01101101;
   assign rom_data[9195]=8'b01010010;
   assign rom_data[9196]=8'b01101101;
   assign rom_data[9197]=8'b01010001;
   assign rom_data[9198]=8'b01101101;
   assign rom_data[9199]=8'b01010000;
   assign rom_data[9200]=8'b01101101;
   assign rom_data[9201]=8'b01001110;
   assign rom_data[9202]=8'b01101101;
   assign rom_data[9203]=8'b01001101;
   assign rom_data[9204]=8'b01101101;
   assign rom_data[9205]=8'b01001100;
   assign rom_data[9206]=8'b01101101;
   assign rom_data[9207]=8'b01001010;
   assign rom_data[9208]=8'b01101101;
   assign rom_data[9209]=8'b01001001;
   assign rom_data[9210]=8'b01101101;
   assign rom_data[9211]=8'b01001000;
   assign rom_data[9212]=8'b01101101;
   assign rom_data[9213]=8'b01000110;
   assign rom_data[9214]=8'b01101101;
   assign rom_data[9215]=8'b01000101;
   assign rom_data[9216]=8'b01101101;
   assign rom_data[9217]=8'b01000100;
   assign rom_data[9218]=8'b01101101;
   assign rom_data[9219]=8'b01000010;
   assign rom_data[9220]=8'b01101100;
   assign rom_data[9221]=8'b01000001;
   assign rom_data[9222]=8'b01101100;
   assign rom_data[9223]=8'b01000000;
   assign rom_data[9224]=8'b01101100;
   assign rom_data[9225]=8'b00111110;
   assign rom_data[9226]=8'b01101100;
   assign rom_data[9227]=8'b00111101;
   assign rom_data[9228]=8'b01101100;
   assign rom_data[9229]=8'b00111100;
   assign rom_data[9230]=8'b01101100;
   assign rom_data[9231]=8'b00111011;
   assign rom_data[9232]=8'b01101100;
   assign rom_data[9233]=8'b00111010;
   assign rom_data[9234]=8'b01101100;
   assign rom_data[9235]=8'b00111001;
   assign rom_data[9236]=8'b01101100;
   assign rom_data[9237]=8'b00110111;
   assign rom_data[9238]=8'b01101100;
   assign rom_data[9239]=8'b00110110;
   assign rom_data[9240]=8'b01101100;
   assign rom_data[9241]=8'b00110101;
   assign rom_data[9242]=8'b01101100;
   assign rom_data[9243]=8'b00110100;
   assign rom_data[9244]=8'b01101100;
   assign rom_data[9245]=8'b00110011;
   assign rom_data[9246]=8'b01101100;
   assign rom_data[9247]=8'b00110011;
   assign rom_data[9248]=8'b01101100;
   assign rom_data[9249]=8'b00110010;
   assign rom_data[9250]=8'b01101100;
   assign rom_data[9251]=8'b00110001;
   assign rom_data[9252]=8'b01101100;
   assign rom_data[9253]=8'b00110000;
   assign rom_data[9254]=8'b01101100;
   assign rom_data[9255]=8'b00101111;
   assign rom_data[9256]=8'b01101100;
   assign rom_data[9257]=8'b00101111;
   assign rom_data[9258]=8'b01101100;
   assign rom_data[9259]=8'b00101110;
   assign rom_data[9260]=8'b01101100;
   assign rom_data[9261]=8'b00101110;
   assign rom_data[9262]=8'b01101100;
   assign rom_data[9263]=8'b00101101;
   assign rom_data[9264]=8'b01101100;
   assign rom_data[9265]=8'b00101101;
   assign rom_data[9266]=8'b01101100;
   assign rom_data[9267]=8'b00101100;
   assign rom_data[9268]=8'b01101100;
   assign rom_data[9269]=8'b00101100;
   assign rom_data[9270]=8'b01101100;
   assign rom_data[9271]=8'b00101100;
   assign rom_data[9272]=8'b01101100;
   assign rom_data[9273]=8'b00101100;
   assign rom_data[9274]=8'b01101100;
   assign rom_data[9275]=8'b00101100;
   assign rom_data[9276]=8'b01101100;
   assign rom_data[9277]=8'b00101100;
   assign rom_data[9278]=8'b01101100;
   assign rom_data[9279]=8'b00101100;
   assign rom_data[9280]=8'b01101100;
   assign rom_data[9281]=8'b00101101;
   assign rom_data[9282]=8'b01101100;
   assign rom_data[9283]=8'b00101101;
   assign rom_data[9284]=8'b01101100;
   assign rom_data[9285]=8'b00101101;
   assign rom_data[9286]=8'b01101011;
   assign rom_data[9287]=8'b00101110;
   assign rom_data[9288]=8'b01101011;
   assign rom_data[9289]=8'b00101111;
   assign rom_data[9290]=8'b01101011;
   assign rom_data[9291]=8'b00101111;
   assign rom_data[9292]=8'b01101011;
   assign rom_data[9293]=8'b00110000;
   assign rom_data[9294]=8'b01101011;
   assign rom_data[9295]=8'b00110001;
   assign rom_data[9296]=8'b01101011;
   assign rom_data[9297]=8'b00110001;
   assign rom_data[9298]=8'b01101011;
   assign rom_data[9299]=8'b00110010;
   assign rom_data[9300]=8'b01101011;
   assign rom_data[9301]=8'b00110011;
   assign rom_data[9302]=8'b01101011;
   assign rom_data[9303]=8'b00110100;
   assign rom_data[9304]=8'b01101011;
   assign rom_data[9305]=8'b00110101;
   assign rom_data[9306]=8'b01101011;
   assign rom_data[9307]=8'b00110110;
   assign rom_data[9308]=8'b01101011;
   assign rom_data[9309]=8'b00110111;
   assign rom_data[9310]=8'b01101011;
   assign rom_data[9311]=8'b00111000;
   assign rom_data[9312]=8'b01101011;
   assign rom_data[9313]=8'b00111010;
   assign rom_data[9314]=8'b01101011;
   assign rom_data[9315]=8'b00111011;
   assign rom_data[9316]=8'b01101011;
   assign rom_data[9317]=8'b00111100;
   assign rom_data[9318]=8'b01101011;
   assign rom_data[9319]=8'b00111101;
   assign rom_data[9320]=8'b01101011;
   assign rom_data[9321]=8'b00111110;
   assign rom_data[9322]=8'b01101011;
   assign rom_data[9323]=8'b01000000;
   assign rom_data[9324]=8'b01101011;
   assign rom_data[9325]=8'b01000001;
   assign rom_data[9326]=8'b01101011;
   assign rom_data[9327]=8'b01000010;
   assign rom_data[9328]=8'b01101011;
   assign rom_data[9329]=8'b01000100;
   assign rom_data[9330]=8'b01101011;
   assign rom_data[9331]=8'b01000101;
   assign rom_data[9332]=8'b01101011;
   assign rom_data[9333]=8'b01000110;
   assign rom_data[9334]=8'b01101011;
   assign rom_data[9335]=8'b01001000;
   assign rom_data[9336]=8'b01101011;
   assign rom_data[9337]=8'b01001001;
   assign rom_data[9338]=8'b01101011;
   assign rom_data[9339]=8'b01001010;
   assign rom_data[9340]=8'b01101011;
   assign rom_data[9341]=8'b01001100;
   assign rom_data[9342]=8'b01101011;
   assign rom_data[9343]=8'b01001101;
   assign rom_data[9344]=8'b01101011;
   assign rom_data[9345]=8'b01001110;
   assign rom_data[9346]=8'b01101011;
   assign rom_data[9347]=8'b01010000;
   assign rom_data[9348]=8'b01101011;
   assign rom_data[9349]=8'b01010001;
   assign rom_data[9350]=8'b01101011;
   assign rom_data[9351]=8'b01010011;
   assign rom_data[9352]=8'b01101011;
   assign rom_data[9353]=8'b01010100;
   assign rom_data[9354]=8'b01101011;
   assign rom_data[9355]=8'b01010101;
   assign rom_data[9356]=8'b01101011;
   assign rom_data[9357]=8'b01010111;
   assign rom_data[9358]=8'b01101011;
   assign rom_data[9359]=8'b01011000;
   assign rom_data[9360]=8'b01101011;
   assign rom_data[9361]=8'b01011010;
   assign rom_data[9362]=8'b01101011;
   assign rom_data[9363]=8'b01011011;
   assign rom_data[9364]=8'b01101011;
   assign rom_data[9365]=8'b01011100;
   assign rom_data[9366]=8'b01101010;
   assign rom_data[9367]=8'b01011110;
   assign rom_data[9368]=8'b01101010;
   assign rom_data[9369]=8'b01011111;
   assign rom_data[9370]=8'b01101010;
   assign rom_data[9371]=8'b01100001;
   assign rom_data[9372]=8'b01101010;
   assign rom_data[9373]=8'b01100010;
   assign rom_data[9374]=8'b01101010;
   assign rom_data[9375]=8'b01100011;
   assign rom_data[9376]=8'b01101010;
   assign rom_data[9377]=8'b01100101;
   assign rom_data[9378]=8'b01101010;
   assign rom_data[9379]=8'b01100110;
   assign rom_data[9380]=8'b01101010;
   assign rom_data[9381]=8'b01101000;
   assign rom_data[9382]=8'b01101010;
   assign rom_data[9383]=8'b01101001;
   assign rom_data[9384]=8'b01101010;
   assign rom_data[9385]=8'b01101010;
   assign rom_data[9386]=8'b01101010;
   assign rom_data[9387]=8'b01101100;
   assign rom_data[9388]=8'b01101010;
   assign rom_data[9389]=8'b01101101;
   assign rom_data[9390]=8'b01101010;
   assign rom_data[9391]=8'b01101110;
   assign rom_data[9392]=8'b01101010;
   assign rom_data[9393]=8'b01110000;
   assign rom_data[9394]=8'b01101010;
   assign rom_data[9395]=8'b01110001;
   assign rom_data[9396]=8'b01101010;
   assign rom_data[9397]=8'b01110010;
   assign rom_data[9398]=8'b01101010;
   assign rom_data[9399]=8'b01110100;
   assign rom_data[9400]=8'b01101010;
   assign rom_data[9401]=8'b01110101;
   assign rom_data[9402]=8'b01101010;
   assign rom_data[9403]=8'b01110110;
   assign rom_data[9404]=8'b01101010;
   assign rom_data[9405]=8'b01110111;
   assign rom_data[9406]=8'b01101010;
   assign rom_data[9407]=8'b01111001;
   assign rom_data[9408]=8'b01101010;
   assign rom_data[9409]=8'b01111010;
   assign rom_data[9410]=8'b01101010;
   assign rom_data[9411]=8'b01111011;
   assign rom_data[9412]=8'b01101010;
   assign rom_data[9413]=8'b01111100;
   assign rom_data[9414]=8'b01101010;
   assign rom_data[9415]=8'b01111101;
   assign rom_data[9416]=8'b01101010;
   assign rom_data[9417]=8'b01111110;
   assign rom_data[9418]=8'b01101010;
   assign rom_data[9419]=8'b01111111;
   assign rom_data[9420]=8'b01101010;
   assign rom_data[9421]=8'b10000000;
   assign rom_data[9422]=8'b01101010;
   assign rom_data[9423]=8'b10000001;
   assign rom_data[9424]=8'b01101010;
   assign rom_data[9425]=8'b10000010;
   assign rom_data[9426]=8'b01101010;
   assign rom_data[9427]=8'b10000011;
   assign rom_data[9428]=8'b01101010;
   assign rom_data[9429]=8'b10000100;
   assign rom_data[9430]=8'b01101010;
   assign rom_data[9431]=8'b10000101;
   assign rom_data[9432]=8'b01101010;
   assign rom_data[9433]=8'b10000110;
   assign rom_data[9434]=8'b01101010;
   assign rom_data[9435]=8'b10000110;
   assign rom_data[9436]=8'b01101010;
   assign rom_data[9437]=8'b10000111;
   assign rom_data[9438]=8'b01101010;
   assign rom_data[9439]=8'b10001000;
   assign rom_data[9440]=8'b01101010;
   assign rom_data[9441]=8'b10001000;
   assign rom_data[9442]=8'b01101001;
   assign rom_data[9443]=8'b10001001;
   assign rom_data[9444]=8'b01101001;
   assign rom_data[9445]=8'b10001001;
   assign rom_data[9446]=8'b01101001;
   assign rom_data[9447]=8'b10001001;
   assign rom_data[9448]=8'b01101001;
   assign rom_data[9449]=8'b10001010;
   assign rom_data[9450]=8'b01101001;
   assign rom_data[9451]=8'b10001010;
   assign rom_data[9452]=8'b01101001;
   assign rom_data[9453]=8'b10001010;
   assign rom_data[9454]=8'b01101001;
   assign rom_data[9455]=8'b10001010;
   assign rom_data[9456]=8'b01101001;
   assign rom_data[9457]=8'b10001010;
   assign rom_data[9458]=8'b01101001;
   assign rom_data[9459]=8'b10001001;
   assign rom_data[9460]=8'b01101001;
   assign rom_data[9461]=8'b10001001;
   assign rom_data[9462]=8'b01101001;
   assign rom_data[9463]=8'b10001001;
   assign rom_data[9464]=8'b01101001;
   assign rom_data[9465]=8'b10001000;
   assign rom_data[9466]=8'b01101001;
   assign rom_data[9467]=8'b10001000;
   assign rom_data[9468]=8'b01101001;
   assign rom_data[9469]=8'b10000111;
   assign rom_data[9470]=8'b01101001;
   assign rom_data[9471]=8'b10000111;
   assign rom_data[9472]=8'b01101001;
   assign rom_data[9473]=8'b10000110;
   assign rom_data[9474]=8'b01101001;
   assign rom_data[9475]=8'b10000101;
   assign rom_data[9476]=8'b01101001;
   assign rom_data[9477]=8'b10000100;
   assign rom_data[9478]=8'b01101001;
   assign rom_data[9479]=8'b10000011;
   assign rom_data[9480]=8'b01101001;
   assign rom_data[9481]=8'b10000011;
   assign rom_data[9482]=8'b01101001;
   assign rom_data[9483]=8'b10000010;
   assign rom_data[9484]=8'b01101001;
   assign rom_data[9485]=8'b10000001;
   assign rom_data[9486]=8'b01101001;
   assign rom_data[9487]=8'b10000000;
   assign rom_data[9488]=8'b01101001;
   assign rom_data[9489]=8'b01111110;
   assign rom_data[9490]=8'b01101001;
   assign rom_data[9491]=8'b01111101;
   assign rom_data[9492]=8'b01101001;
   assign rom_data[9493]=8'b01111100;
   assign rom_data[9494]=8'b01101001;
   assign rom_data[9495]=8'b01111011;
   assign rom_data[9496]=8'b01101001;
   assign rom_data[9497]=8'b01111010;
   assign rom_data[9498]=8'b01101001;
   assign rom_data[9499]=8'b01111001;
   assign rom_data[9500]=8'b01101001;
   assign rom_data[9501]=8'b01110111;
   assign rom_data[9502]=8'b01101001;
   assign rom_data[9503]=8'b01110110;
   assign rom_data[9504]=8'b01101001;
   assign rom_data[9505]=8'b01110101;
   assign rom_data[9506]=8'b01101001;
   assign rom_data[9507]=8'b01110100;
   assign rom_data[9508]=8'b01101001;
   assign rom_data[9509]=8'b01110010;
   assign rom_data[9510]=8'b01101000;
   assign rom_data[9511]=8'b01110001;
   assign rom_data[9512]=8'b01101000;
   assign rom_data[9513]=8'b01110000;
   assign rom_data[9514]=8'b01101000;
   assign rom_data[9515]=8'b01101110;
   assign rom_data[9516]=8'b01101000;
   assign rom_data[9517]=8'b01101101;
   assign rom_data[9518]=8'b01101000;
   assign rom_data[9519]=8'b01101100;
   assign rom_data[9520]=8'b01101000;
   assign rom_data[9521]=8'b01101010;
   assign rom_data[9522]=8'b01101000;
   assign rom_data[9523]=8'b01101001;
   assign rom_data[9524]=8'b01101000;
   assign rom_data[9525]=8'b01100111;
   assign rom_data[9526]=8'b01101000;
   assign rom_data[9527]=8'b01100110;
   assign rom_data[9528]=8'b01101000;
   assign rom_data[9529]=8'b01100101;
   assign rom_data[9530]=8'b01101000;
   assign rom_data[9531]=8'b01100011;
   assign rom_data[9532]=8'b01101000;
   assign rom_data[9533]=8'b01100010;
   assign rom_data[9534]=8'b01101000;
   assign rom_data[9535]=8'b01100000;
   assign rom_data[9536]=8'b01101000;
   assign rom_data[9537]=8'b01011111;
   assign rom_data[9538]=8'b01101000;
   assign rom_data[9539]=8'b01011110;
   assign rom_data[9540]=8'b01101000;
   assign rom_data[9541]=8'b01011100;
   assign rom_data[9542]=8'b01101000;
   assign rom_data[9543]=8'b01011011;
   assign rom_data[9544]=8'b01101000;
   assign rom_data[9545]=8'b01011001;
   assign rom_data[9546]=8'b01101000;
   assign rom_data[9547]=8'b01011000;
   assign rom_data[9548]=8'b01101000;
   assign rom_data[9549]=8'b01010111;
   assign rom_data[9550]=8'b01101000;
   assign rom_data[9551]=8'b01010101;
   assign rom_data[9552]=8'b01101000;
   assign rom_data[9553]=8'b01010100;
   assign rom_data[9554]=8'b01101000;
   assign rom_data[9555]=8'b01010010;
   assign rom_data[9556]=8'b01101000;
   assign rom_data[9557]=8'b01010001;
   assign rom_data[9558]=8'b01101000;
   assign rom_data[9559]=8'b01010000;
   assign rom_data[9560]=8'b01101000;
   assign rom_data[9561]=8'b01001110;
   assign rom_data[9562]=8'b01101000;
   assign rom_data[9563]=8'b01001101;
   assign rom_data[9564]=8'b01101000;
   assign rom_data[9565]=8'b01001100;
   assign rom_data[9566]=8'b01101000;
   assign rom_data[9567]=8'b01001010;
   assign rom_data[9568]=8'b01101000;
   assign rom_data[9569]=8'b01001001;
   assign rom_data[9570]=8'b01101000;
   assign rom_data[9571]=8'b01001000;
   assign rom_data[9572]=8'b01101000;
   assign rom_data[9573]=8'b01000110;
   assign rom_data[9574]=8'b01101000;
   assign rom_data[9575]=8'b01000101;
   assign rom_data[9576]=8'b01101000;
   assign rom_data[9577]=8'b01000100;
   assign rom_data[9578]=8'b01101000;
   assign rom_data[9579]=8'b01000010;
   assign rom_data[9580]=8'b01101000;
   assign rom_data[9581]=8'b01000001;
   assign rom_data[9582]=8'b01101000;
   assign rom_data[9583]=8'b01000000;
   assign rom_data[9584]=8'b01101000;
   assign rom_data[9585]=8'b00111110;
   assign rom_data[9586]=8'b01101000;
   assign rom_data[9587]=8'b00111101;
   assign rom_data[9588]=8'b01101000;
   assign rom_data[9589]=8'b00111100;
   assign rom_data[9590]=8'b01101000;
   assign rom_data[9591]=8'b00111011;
   assign rom_data[9592]=8'b01101000;
   assign rom_data[9593]=8'b00111010;
   assign rom_data[9594]=8'b01100111;
   assign rom_data[9595]=8'b00111001;
   assign rom_data[9596]=8'b01100111;
   assign rom_data[9597]=8'b00110111;
   assign rom_data[9598]=8'b01100111;
   assign rom_data[9599]=8'b00110110;
   assign rom_data[9600]=8'b01100111;
   assign rom_data[9601]=8'b00110101;
   assign rom_data[9602]=8'b01100111;
   assign rom_data[9603]=8'b00110100;
   assign rom_data[9604]=8'b01100111;
   assign rom_data[9605]=8'b00110011;
   assign rom_data[9606]=8'b01100111;
   assign rom_data[9607]=8'b00110011;
   assign rom_data[9608]=8'b01100111;
   assign rom_data[9609]=8'b00110010;
   assign rom_data[9610]=8'b01100111;
   assign rom_data[9611]=8'b00110001;
   assign rom_data[9612]=8'b01100111;
   assign rom_data[9613]=8'b00110000;
   assign rom_data[9614]=8'b01100111;
   assign rom_data[9615]=8'b00101111;
   assign rom_data[9616]=8'b01100111;
   assign rom_data[9617]=8'b00101111;
   assign rom_data[9618]=8'b01100111;
   assign rom_data[9619]=8'b00101110;
   assign rom_data[9620]=8'b01100111;
   assign rom_data[9621]=8'b00101110;
   assign rom_data[9622]=8'b01100111;
   assign rom_data[9623]=8'b00101101;
   assign rom_data[9624]=8'b01100111;
   assign rom_data[9625]=8'b00101101;
   assign rom_data[9626]=8'b01100111;
   assign rom_data[9627]=8'b00101100;
   assign rom_data[9628]=8'b01100111;
   assign rom_data[9629]=8'b00101100;
   assign rom_data[9630]=8'b01100111;
   assign rom_data[9631]=8'b00101100;
   assign rom_data[9632]=8'b01100111;
   assign rom_data[9633]=8'b00101100;
   assign rom_data[9634]=8'b01100111;
   assign rom_data[9635]=8'b00101100;
   assign rom_data[9636]=8'b01100111;
   assign rom_data[9637]=8'b00101100;
   assign rom_data[9638]=8'b01100111;
   assign rom_data[9639]=8'b00101100;
   assign rom_data[9640]=8'b01100111;
   assign rom_data[9641]=8'b00101101;
   assign rom_data[9642]=8'b01100111;
   assign rom_data[9643]=8'b00101101;
   assign rom_data[9644]=8'b01100111;
   assign rom_data[9645]=8'b00101101;
   assign rom_data[9646]=8'b01100111;
   assign rom_data[9647]=8'b00101110;
   assign rom_data[9648]=8'b01100111;
   assign rom_data[9649]=8'b00101111;
   assign rom_data[9650]=8'b01100111;
   assign rom_data[9651]=8'b00101111;
   assign rom_data[9652]=8'b01100111;
   assign rom_data[9653]=8'b00110000;
   assign rom_data[9654]=8'b01100111;
   assign rom_data[9655]=8'b00110001;
   assign rom_data[9656]=8'b01100111;
   assign rom_data[9657]=8'b00110001;
   assign rom_data[9658]=8'b01100111;
   assign rom_data[9659]=8'b00110010;
   assign rom_data[9660]=8'b01100110;
   assign rom_data[9661]=8'b00110011;
   assign rom_data[9662]=8'b01100110;
   assign rom_data[9663]=8'b00110100;
   assign rom_data[9664]=8'b01100110;
   assign rom_data[9665]=8'b00110101;
   assign rom_data[9666]=8'b01100110;
   assign rom_data[9667]=8'b00110110;
   assign rom_data[9668]=8'b01100110;
   assign rom_data[9669]=8'b00110111;
   assign rom_data[9670]=8'b01100110;
   assign rom_data[9671]=8'b00111000;
   assign rom_data[9672]=8'b01100110;
   assign rom_data[9673]=8'b00111010;
   assign rom_data[9674]=8'b01100110;
   assign rom_data[9675]=8'b00111011;
   assign rom_data[9676]=8'b01100110;
   assign rom_data[9677]=8'b00111100;
   assign rom_data[9678]=8'b01100110;
   assign rom_data[9679]=8'b00111101;
   assign rom_data[9680]=8'b01100110;
   assign rom_data[9681]=8'b00111110;
   assign rom_data[9682]=8'b01100110;
   assign rom_data[9683]=8'b01000000;
   assign rom_data[9684]=8'b01100110;
   assign rom_data[9685]=8'b01000001;
   assign rom_data[9686]=8'b01100110;
   assign rom_data[9687]=8'b01000010;
   assign rom_data[9688]=8'b01100110;
   assign rom_data[9689]=8'b01000100;
   assign rom_data[9690]=8'b01100110;
   assign rom_data[9691]=8'b01000101;
   assign rom_data[9692]=8'b01100110;
   assign rom_data[9693]=8'b01000110;
   assign rom_data[9694]=8'b01100110;
   assign rom_data[9695]=8'b01001000;
   assign rom_data[9696]=8'b01100110;
   assign rom_data[9697]=8'b01001001;
   assign rom_data[9698]=8'b01100110;
   assign rom_data[9699]=8'b01001010;
   assign rom_data[9700]=8'b01100110;
   assign rom_data[9701]=8'b01001100;
   assign rom_data[9702]=8'b01100110;
   assign rom_data[9703]=8'b01001101;
   assign rom_data[9704]=8'b01100110;
   assign rom_data[9705]=8'b01001110;
   assign rom_data[9706]=8'b01100110;
   assign rom_data[9707]=8'b01010000;
   assign rom_data[9708]=8'b01100110;
   assign rom_data[9709]=8'b01010001;
   assign rom_data[9710]=8'b01100110;
   assign rom_data[9711]=8'b01010011;
   assign rom_data[9712]=8'b01100110;
   assign rom_data[9713]=8'b01010100;
   assign rom_data[9714]=8'b01100110;
   assign rom_data[9715]=8'b01010101;
   assign rom_data[9716]=8'b01100110;
   assign rom_data[9717]=8'b01010111;
   assign rom_data[9718]=8'b01100110;
   assign rom_data[9719]=8'b01011000;
   assign rom_data[9720]=8'b01100110;
   assign rom_data[9721]=8'b01011010;
   assign rom_data[9722]=8'b01100110;
   assign rom_data[9723]=8'b01011011;
   assign rom_data[9724]=8'b01100110;
   assign rom_data[9725]=8'b01011100;
   assign rom_data[9726]=8'b01100110;
   assign rom_data[9727]=8'b01011110;
   assign rom_data[9728]=8'b01100110;
   assign rom_data[9729]=8'b01011111;
   assign rom_data[9730]=8'b01100110;
   assign rom_data[9731]=8'b01100001;
   assign rom_data[9732]=8'b01100110;
   assign rom_data[9733]=8'b01100010;
   assign rom_data[9734]=8'b01100110;
   assign rom_data[9735]=8'b01100011;
   assign rom_data[9736]=8'b01100110;
   assign rom_data[9737]=8'b01100101;
   assign rom_data[9738]=8'b01100110;
   assign rom_data[9739]=8'b01100110;
   assign rom_data[9740]=8'b01100110;
   assign rom_data[9741]=8'b01101000;
   assign rom_data[9742]=8'b01100101;
   assign rom_data[9743]=8'b01101001;
   assign rom_data[9744]=8'b01100101;
   assign rom_data[9745]=8'b01101010;
   assign rom_data[9746]=8'b01100101;
   assign rom_data[9747]=8'b01101100;
   assign rom_data[9748]=8'b01100101;
   assign rom_data[9749]=8'b01101101;
   assign rom_data[9750]=8'b01100101;
   assign rom_data[9751]=8'b01101110;
   assign rom_data[9752]=8'b01100101;
   assign rom_data[9753]=8'b01110000;
   assign rom_data[9754]=8'b01100101;
   assign rom_data[9755]=8'b01110001;
   assign rom_data[9756]=8'b01100101;
   assign rom_data[9757]=8'b01110010;
   assign rom_data[9758]=8'b01100101;
   assign rom_data[9759]=8'b01110100;
   assign rom_data[9760]=8'b01100101;
   assign rom_data[9761]=8'b01110101;
   assign rom_data[9762]=8'b01100101;
   assign rom_data[9763]=8'b01110110;
   assign rom_data[9764]=8'b01100101;
   assign rom_data[9765]=8'b01110111;
   assign rom_data[9766]=8'b01100101;
   assign rom_data[9767]=8'b01111001;
   assign rom_data[9768]=8'b01100101;
   assign rom_data[9769]=8'b01111010;
   assign rom_data[9770]=8'b01100101;
   assign rom_data[9771]=8'b01111011;
   assign rom_data[9772]=8'b01100101;
   assign rom_data[9773]=8'b01111100;
   assign rom_data[9774]=8'b01100101;
   assign rom_data[9775]=8'b01111101;
   assign rom_data[9776]=8'b01100101;
   assign rom_data[9777]=8'b01111110;
   assign rom_data[9778]=8'b01100101;
   assign rom_data[9779]=8'b01111111;
   assign rom_data[9780]=8'b01100101;
   assign rom_data[9781]=8'b10000000;
   assign rom_data[9782]=8'b01100101;
   assign rom_data[9783]=8'b10000001;
   assign rom_data[9784]=8'b01100101;
   assign rom_data[9785]=8'b10000010;
   assign rom_data[9786]=8'b01100101;
   assign rom_data[9787]=8'b10000011;
   assign rom_data[9788]=8'b01100101;
   assign rom_data[9789]=8'b10000100;
   assign rom_data[9790]=8'b01100101;
   assign rom_data[9791]=8'b10000101;
   assign rom_data[9792]=8'b01100101;
   assign rom_data[9793]=8'b10000110;
   assign rom_data[9794]=8'b01100101;
   assign rom_data[9795]=8'b10000110;
   assign rom_data[9796]=8'b01100101;
   assign rom_data[9797]=8'b10000111;
   assign rom_data[9798]=8'b01100101;
   assign rom_data[9799]=8'b10001000;
   assign rom_data[9800]=8'b01100101;
   assign rom_data[9801]=8'b10001000;
   assign rom_data[9802]=8'b01100101;
   assign rom_data[9803]=8'b10001001;
   assign rom_data[9804]=8'b01100101;
   assign rom_data[9805]=8'b10001001;
   assign rom_data[9806]=8'b01100101;
   assign rom_data[9807]=8'b10001001;
   assign rom_data[9808]=8'b01100101;
   assign rom_data[9809]=8'b10001010;
   assign rom_data[9810]=8'b01100101;
   assign rom_data[9811]=8'b10001010;
   assign rom_data[9812]=8'b01100100;
   assign rom_data[9813]=8'b10001010;
   assign rom_data[9814]=8'b01100100;
   assign rom_data[9815]=8'b10001010;
   assign rom_data[9816]=8'b01100100;
   assign rom_data[9817]=8'b10001010;
   assign rom_data[9818]=8'b01100100;
   assign rom_data[9819]=8'b10001001;
   assign rom_data[9820]=8'b01100100;
   assign rom_data[9821]=8'b10001001;
   assign rom_data[9822]=8'b01100100;
   assign rom_data[9823]=8'b10001001;
   assign rom_data[9824]=8'b01100100;
   assign rom_data[9825]=8'b10001000;
   assign rom_data[9826]=8'b01100100;
   assign rom_data[9827]=8'b10001000;
   assign rom_data[9828]=8'b01100100;
   assign rom_data[9829]=8'b10000111;
   assign rom_data[9830]=8'b01100100;
   assign rom_data[9831]=8'b10000111;
   assign rom_data[9832]=8'b01100100;
   assign rom_data[9833]=8'b10000110;
   assign rom_data[9834]=8'b01100100;
   assign rom_data[9835]=8'b10000101;
   assign rom_data[9836]=8'b01100100;
   assign rom_data[9837]=8'b10000100;
   assign rom_data[9838]=8'b01100100;
   assign rom_data[9839]=8'b10000011;
   assign rom_data[9840]=8'b01100100;
   assign rom_data[9841]=8'b10000011;
   assign rom_data[9842]=8'b01100100;
   assign rom_data[9843]=8'b10000010;
   assign rom_data[9844]=8'b01100100;
   assign rom_data[9845]=8'b10000001;
   assign rom_data[9846]=8'b01100100;
   assign rom_data[9847]=8'b10000000;
   assign rom_data[9848]=8'b01100100;
   assign rom_data[9849]=8'b01111110;
   assign rom_data[9850]=8'b01100100;
   assign rom_data[9851]=8'b01111101;
   assign rom_data[9852]=8'b01100100;
   assign rom_data[9853]=8'b01111100;
   assign rom_data[9854]=8'b01100100;
   assign rom_data[9855]=8'b01111011;
   assign rom_data[9856]=8'b01100100;
   assign rom_data[9857]=8'b01111010;
   assign rom_data[9858]=8'b01100100;
   assign rom_data[9859]=8'b01111001;
   assign rom_data[9860]=8'b01100100;
   assign rom_data[9861]=8'b01110111;
   assign rom_data[9862]=8'b01100100;
   assign rom_data[9863]=8'b01110110;
   assign rom_data[9864]=8'b01100100;
   assign rom_data[9865]=8'b01110101;
   assign rom_data[9866]=8'b01100100;
   assign rom_data[9867]=8'b01110100;
   assign rom_data[9868]=8'b01100100;
   assign rom_data[9869]=8'b01110010;
   assign rom_data[9870]=8'b01100100;
   assign rom_data[9871]=8'b01110001;
   assign rom_data[9872]=8'b01100100;
   assign rom_data[9873]=8'b01110000;
   assign rom_data[9874]=8'b01100100;
   assign rom_data[9875]=8'b01101110;
   assign rom_data[9876]=8'b01100100;
   assign rom_data[9877]=8'b01101101;
   assign rom_data[9878]=8'b01100100;
   assign rom_data[9879]=8'b01101100;
   assign rom_data[9880]=8'b01100100;
   assign rom_data[9881]=8'b01101010;
   assign rom_data[9882]=8'b01100100;
   assign rom_data[9883]=8'b01101001;
   assign rom_data[9884]=8'b01100100;
   assign rom_data[9885]=8'b01100111;
   assign rom_data[9886]=8'b01100011;
   assign rom_data[9887]=8'b01100110;
   assign rom_data[9888]=8'b01100011;
   assign rom_data[9889]=8'b01100101;
   assign rom_data[9890]=8'b01100011;
   assign rom_data[9891]=8'b01100011;
   assign rom_data[9892]=8'b01100011;
   assign rom_data[9893]=8'b01100010;
   assign rom_data[9894]=8'b01100011;
   assign rom_data[9895]=8'b01100000;
   assign rom_data[9896]=8'b01100011;
   assign rom_data[9897]=8'b01011111;
   assign rom_data[9898]=8'b01100011;
   assign rom_data[9899]=8'b01011110;
   assign rom_data[9900]=8'b01100011;
   assign rom_data[9901]=8'b01011100;
   assign rom_data[9902]=8'b01100011;
   assign rom_data[9903]=8'b01011011;
   assign rom_data[9904]=8'b01100011;
   assign rom_data[9905]=8'b01011001;
   assign rom_data[9906]=8'b01100011;
   assign rom_data[9907]=8'b01011000;
   assign rom_data[9908]=8'b01100011;
   assign rom_data[9909]=8'b01010111;
   assign rom_data[9910]=8'b01100011;
   assign rom_data[9911]=8'b01010101;
   assign rom_data[9912]=8'b01100011;
   assign rom_data[9913]=8'b01010100;
   assign rom_data[9914]=8'b01100011;
   assign rom_data[9915]=8'b01010010;
   assign rom_data[9916]=8'b01100011;
   assign rom_data[9917]=8'b01010001;
   assign rom_data[9918]=8'b01100011;
   assign rom_data[9919]=8'b01010000;
   assign rom_data[9920]=8'b01100011;
   assign rom_data[9921]=8'b01001110;
   assign rom_data[9922]=8'b01100011;
   assign rom_data[9923]=8'b01001101;
   assign rom_data[9924]=8'b01100011;
   assign rom_data[9925]=8'b01001100;
   assign rom_data[9926]=8'b01100011;
   assign rom_data[9927]=8'b01001010;
   assign rom_data[9928]=8'b01100011;
   assign rom_data[9929]=8'b01001001;
   assign rom_data[9930]=8'b01100011;
   assign rom_data[9931]=8'b01000111;
   assign rom_data[9932]=8'b01100011;
   assign rom_data[9933]=8'b01000110;
   assign rom_data[9934]=8'b01100011;
   assign rom_data[9935]=8'b01000101;
   assign rom_data[9936]=8'b01100011;
   assign rom_data[9937]=8'b01000100;
   assign rom_data[9938]=8'b01100011;
   assign rom_data[9939]=8'b01000010;
   assign rom_data[9940]=8'b01100011;
   assign rom_data[9941]=8'b01000001;
   assign rom_data[9942]=8'b01100011;
   assign rom_data[9943]=8'b01000000;
   assign rom_data[9944]=8'b01100011;
   assign rom_data[9945]=8'b00111110;
   assign rom_data[9946]=8'b01100011;
   assign rom_data[9947]=8'b00111101;
   assign rom_data[9948]=8'b01100011;
   assign rom_data[9949]=8'b00111100;
   assign rom_data[9950]=8'b01100011;
   assign rom_data[9951]=8'b00111011;
   assign rom_data[9952]=8'b01100011;
   assign rom_data[9953]=8'b00111010;
   assign rom_data[9954]=8'b01100011;
   assign rom_data[9955]=8'b00111001;
   assign rom_data[9956]=8'b01100011;
   assign rom_data[9957]=8'b00110111;
   assign rom_data[9958]=8'b01100011;
   assign rom_data[9959]=8'b00110110;
   assign rom_data[9960]=8'b01100011;
   assign rom_data[9961]=8'b00110101;
   assign rom_data[9962]=8'b01100011;
   assign rom_data[9963]=8'b00110100;
   assign rom_data[9964]=8'b01100011;
   assign rom_data[9965]=8'b00110011;
   assign rom_data[9966]=8'b01100011;
   assign rom_data[9967]=8'b00110011;
   assign rom_data[9968]=8'b01100010;
   assign rom_data[9969]=8'b00110010;
   assign rom_data[9970]=8'b01100010;
   assign rom_data[9971]=8'b00110001;
   assign rom_data[9972]=8'b01100010;
   assign rom_data[9973]=8'b00110000;
   assign rom_data[9974]=8'b01100010;
   assign rom_data[9975]=8'b00101111;
   assign rom_data[9976]=8'b01100010;
   assign rom_data[9977]=8'b00101111;
   assign rom_data[9978]=8'b01100010;
   assign rom_data[9979]=8'b00101110;
   assign rom_data[9980]=8'b01100010;
   assign rom_data[9981]=8'b00101110;
   assign rom_data[9982]=8'b01100010;
   assign rom_data[9983]=8'b00101101;
   assign rom_data[9984]=8'b01100010;
   assign rom_data[9985]=8'b00101101;
   assign rom_data[9986]=8'b01100010;
   assign rom_data[9987]=8'b00101100;
   assign rom_data[9988]=8'b01100010;
   assign rom_data[9989]=8'b00101100;
   assign rom_data[9990]=8'b01100010;
   assign rom_data[9991]=8'b00101100;
   assign rom_data[9992]=8'b01100010;
   assign rom_data[9993]=8'b00101100;
   assign rom_data[9994]=8'b01100010;
   assign rom_data[9995]=8'b00101100;
   assign rom_data[9996]=8'b01100010;
   assign rom_data[9997]=8'b00101100;
   assign rom_data[9998]=8'b01100010;
   assign rom_data[9999]=8'b00101100;
   assign rom_data[10000]=8'b01100010;
   assign rom_data[10001]=8'b00101101;
   assign rom_data[10002]=8'b01100010;
   assign rom_data[10003]=8'b00101101;
   assign rom_data[10004]=8'b01100010;
   assign rom_data[10005]=8'b00101101;
   assign rom_data[10006]=8'b01100010;
   assign rom_data[10007]=8'b00101110;
   assign rom_data[10008]=8'b01100010;
   assign rom_data[10009]=8'b00101111;
   assign rom_data[10010]=8'b01100010;
   assign rom_data[10011]=8'b00101111;
   assign rom_data[10012]=8'b01100010;
   assign rom_data[10013]=8'b00110000;
   assign rom_data[10014]=8'b01100010;
   assign rom_data[10015]=8'b00110001;
   assign rom_data[10016]=8'b01100010;
   assign rom_data[10017]=8'b00110001;
   assign rom_data[10018]=8'b01100010;
   assign rom_data[10019]=8'b00110010;
   assign rom_data[10020]=8'b01100010;
   assign rom_data[10021]=8'b00110011;
   assign rom_data[10022]=8'b01100010;
   assign rom_data[10023]=8'b00110100;
   assign rom_data[10024]=8'b01100010;
   assign rom_data[10025]=8'b00110101;
   assign rom_data[10026]=8'b01100010;
   assign rom_data[10027]=8'b00110110;
   assign rom_data[10028]=8'b01100010;
   assign rom_data[10029]=8'b00110111;
   assign rom_data[10030]=8'b01100010;
   assign rom_data[10031]=8'b00111000;
   assign rom_data[10032]=8'b01100010;
   assign rom_data[10033]=8'b00111010;
   assign rom_data[10034]=8'b01100001;
   assign rom_data[10035]=8'b00111011;
   assign rom_data[10036]=8'b01100001;
   assign rom_data[10037]=8'b00111100;
   assign rom_data[10038]=8'b01100001;
   assign rom_data[10039]=8'b00111101;
   assign rom_data[10040]=8'b01100001;
   assign rom_data[10041]=8'b00111110;
   assign rom_data[10042]=8'b01100001;
   assign rom_data[10043]=8'b01000000;
   assign rom_data[10044]=8'b01100001;
   assign rom_data[10045]=8'b01000001;
   assign rom_data[10046]=8'b01100001;
   assign rom_data[10047]=8'b01000010;
   assign rom_data[10048]=8'b01100001;
   assign rom_data[10049]=8'b01000100;
   assign rom_data[10050]=8'b01100001;
   assign rom_data[10051]=8'b01000101;
   assign rom_data[10052]=8'b01100001;
   assign rom_data[10053]=8'b01000110;
   assign rom_data[10054]=8'b01100001;
   assign rom_data[10055]=8'b01001000;
   assign rom_data[10056]=8'b01100001;
   assign rom_data[10057]=8'b01001001;
   assign rom_data[10058]=8'b01100001;
   assign rom_data[10059]=8'b01001010;
   assign rom_data[10060]=8'b01100001;
   assign rom_data[10061]=8'b01001100;
   assign rom_data[10062]=8'b01100001;
   assign rom_data[10063]=8'b01001101;
   assign rom_data[10064]=8'b01100001;
   assign rom_data[10065]=8'b01001110;
   assign rom_data[10066]=8'b01100001;
   assign rom_data[10067]=8'b01010000;
   assign rom_data[10068]=8'b01100001;
   assign rom_data[10069]=8'b01010001;
   assign rom_data[10070]=8'b01100001;
   assign rom_data[10071]=8'b01010011;
   assign rom_data[10072]=8'b01100001;
   assign rom_data[10073]=8'b01010100;
   assign rom_data[10074]=8'b01100001;
   assign rom_data[10075]=8'b01010101;
   assign rom_data[10076]=8'b01100001;
   assign rom_data[10077]=8'b01010111;
   assign rom_data[10078]=8'b01100001;
   assign rom_data[10079]=8'b01011000;
   assign rom_data[10080]=8'b01100001;
   assign rom_data[10081]=8'b01011010;
   assign rom_data[10082]=8'b01100001;
   assign rom_data[10083]=8'b01011011;
   assign rom_data[10084]=8'b01100001;
   assign rom_data[10085]=8'b01011100;
   assign rom_data[10086]=8'b01100001;
   assign rom_data[10087]=8'b01011110;
   assign rom_data[10088]=8'b01100001;
   assign rom_data[10089]=8'b01011111;
   assign rom_data[10090]=8'b01100001;
   assign rom_data[10091]=8'b01100001;
   assign rom_data[10092]=8'b01100001;
   assign rom_data[10093]=8'b01100010;
   assign rom_data[10094]=8'b01100001;
   assign rom_data[10095]=8'b01100011;
   assign rom_data[10096]=8'b01100001;
   assign rom_data[10097]=8'b01100101;
   assign rom_data[10098]=8'b01100001;
   assign rom_data[10099]=8'b01100110;
   assign rom_data[10100]=8'b01100001;
   assign rom_data[10101]=8'b01101000;
   assign rom_data[10102]=8'b01100001;
   assign rom_data[10103]=8'b01101001;
   assign rom_data[10104]=8'b01100001;
   assign rom_data[10105]=8'b01101010;
   assign rom_data[10106]=8'b01100001;
   assign rom_data[10107]=8'b01101100;
   assign rom_data[10108]=8'b01100001;
   assign rom_data[10109]=8'b01101101;
   assign rom_data[10110]=8'b01100001;
   assign rom_data[10111]=8'b01101110;
   assign rom_data[10112]=8'b01100001;
   assign rom_data[10113]=8'b01110000;
   assign rom_data[10114]=8'b01100001;
   assign rom_data[10115]=8'b01110001;
   assign rom_data[10116]=8'b01100001;
   assign rom_data[10117]=8'b01110010;
   assign rom_data[10118]=8'b01100000;
   assign rom_data[10119]=8'b01110100;
   assign rom_data[10120]=8'b01100000;
   assign rom_data[10121]=8'b01110101;
   assign rom_data[10122]=8'b01100000;
   assign rom_data[10123]=8'b01110110;
   assign rom_data[10124]=8'b01100000;
   assign rom_data[10125]=8'b01110111;
   assign rom_data[10126]=8'b01100000;
   assign rom_data[10127]=8'b01111001;
   assign rom_data[10128]=8'b01100000;
   assign rom_data[10129]=8'b01111010;
   assign rom_data[10130]=8'b01100000;
   assign rom_data[10131]=8'b01111011;
   assign rom_data[10132]=8'b01100000;
   assign rom_data[10133]=8'b01111100;
   assign rom_data[10134]=8'b01100000;
   assign rom_data[10135]=8'b01111101;
   assign rom_data[10136]=8'b01100000;
   assign rom_data[10137]=8'b01111110;
   assign rom_data[10138]=8'b01100000;
   assign rom_data[10139]=8'b01111111;
   assign rom_data[10140]=8'b01100000;
   assign rom_data[10141]=8'b10000000;
   assign rom_data[10142]=8'b01100000;
   assign rom_data[10143]=8'b10000001;
   assign rom_data[10144]=8'b01100000;
   assign rom_data[10145]=8'b10000010;
   assign rom_data[10146]=8'b01100000;
   assign rom_data[10147]=8'b10000011;
   assign rom_data[10148]=8'b01100000;
   assign rom_data[10149]=8'b10000100;
   assign rom_data[10150]=8'b01100000;
   assign rom_data[10151]=8'b10000101;
   assign rom_data[10152]=8'b01100000;
   assign rom_data[10153]=8'b10000110;
   assign rom_data[10154]=8'b01100000;
   assign rom_data[10155]=8'b10000110;
   assign rom_data[10156]=8'b01100000;
   assign rom_data[10157]=8'b10000111;
   assign rom_data[10158]=8'b01100000;
   assign rom_data[10159]=8'b10001000;
   assign rom_data[10160]=8'b01100000;
   assign rom_data[10161]=8'b10001000;
   assign rom_data[10162]=8'b01100000;
   assign rom_data[10163]=8'b10001001;
   assign rom_data[10164]=8'b01100000;
   assign rom_data[10165]=8'b10001001;
   assign rom_data[10166]=8'b01100000;
   assign rom_data[10167]=8'b10001001;
   assign rom_data[10168]=8'b01100000;
   assign rom_data[10169]=8'b10001010;
   assign rom_data[10170]=8'b01100000;
   assign rom_data[10171]=8'b10001010;
   assign rom_data[10172]=8'b01100000;
   assign rom_data[10173]=8'b10001010;
   assign rom_data[10174]=8'b01100000;
   assign rom_data[10175]=8'b10001010;
   assign rom_data[10176]=8'b01100000;
   assign rom_data[10177]=8'b10001010;
   assign rom_data[10178]=8'b01100000;
   assign rom_data[10179]=8'b10001001;
   assign rom_data[10180]=8'b01100000;
   assign rom_data[10181]=8'b10001001;
   assign rom_data[10182]=8'b01100000;
   assign rom_data[10183]=8'b10001001;
   assign rom_data[10184]=8'b01011111;
   assign rom_data[10185]=8'b10001000;
   assign rom_data[10186]=8'b01011111;
   assign rom_data[10187]=8'b10001000;
   assign rom_data[10188]=8'b01011111;
   assign rom_data[10189]=8'b10000111;
   assign rom_data[10190]=8'b01011111;
   assign rom_data[10191]=8'b10000111;
   assign rom_data[10192]=8'b01011111;
   assign rom_data[10193]=8'b10000110;
   assign rom_data[10194]=8'b01011111;
   assign rom_data[10195]=8'b10000101;
   assign rom_data[10196]=8'b01011111;
   assign rom_data[10197]=8'b10000100;
   assign rom_data[10198]=8'b01011111;
   assign rom_data[10199]=8'b10000011;
   assign rom_data[10200]=8'b01011111;
   assign rom_data[10201]=8'b10000011;
   assign rom_data[10202]=8'b01011111;
   assign rom_data[10203]=8'b10000010;
   assign rom_data[10204]=8'b01011111;
   assign rom_data[10205]=8'b10000001;
   assign rom_data[10206]=8'b01011111;
   assign rom_data[10207]=8'b10000000;
   assign rom_data[10208]=8'b01011111;
   assign rom_data[10209]=8'b01111110;
   assign rom_data[10210]=8'b01011111;
   assign rom_data[10211]=8'b01111101;
   assign rom_data[10212]=8'b01011111;
   assign rom_data[10213]=8'b01111100;
   assign rom_data[10214]=8'b01011111;
   assign rom_data[10215]=8'b01111011;
   assign rom_data[10216]=8'b01011111;
   assign rom_data[10217]=8'b01111010;
   assign rom_data[10218]=8'b01011111;
   assign rom_data[10219]=8'b01111001;
   assign rom_data[10220]=8'b01011111;
   assign rom_data[10221]=8'b01110111;
   assign rom_data[10222]=8'b01011111;
   assign rom_data[10223]=8'b01110110;
   assign rom_data[10224]=8'b01011111;
   assign rom_data[10225]=8'b01110101;
   assign rom_data[10226]=8'b01011111;
   assign rom_data[10227]=8'b01110100;
   assign rom_data[10228]=8'b01011111;
   assign rom_data[10229]=8'b01110010;
   assign rom_data[10230]=8'b01011111;
   assign rom_data[10231]=8'b01110001;
   assign rom_data[10232]=8'b01011111;
   assign rom_data[10233]=8'b01110000;
   assign rom_data[10234]=8'b01011111;
   assign rom_data[10235]=8'b01101110;
   assign rom_data[10236]=8'b01011111;
   assign rom_data[10237]=8'b01101101;
   assign rom_data[10238]=8'b01011111;
   assign rom_data[10239]=8'b01101100;
   assign rom_data[10240]=8'b01011111;
   assign rom_data[10241]=8'b01101010;
   assign rom_data[10242]=8'b01011111;
   assign rom_data[10243]=8'b01101001;
   assign rom_data[10244]=8'b01011111;
   assign rom_data[10245]=8'b01100111;
   assign rom_data[10246]=8'b01011111;
   assign rom_data[10247]=8'b01100110;
   assign rom_data[10248]=8'b01011111;
   assign rom_data[10249]=8'b01100101;
   assign rom_data[10250]=8'b01011111;
   assign rom_data[10251]=8'b01100011;
   assign rom_data[10252]=8'b01011111;
   assign rom_data[10253]=8'b01100010;
   assign rom_data[10254]=8'b01011111;
   assign rom_data[10255]=8'b01100000;
   assign rom_data[10256]=8'b01011111;
   assign rom_data[10257]=8'b01011111;
   assign rom_data[10258]=8'b01011111;
   assign rom_data[10259]=8'b01011110;
   assign rom_data[10260]=8'b01011111;
   assign rom_data[10261]=8'b01011100;
   assign rom_data[10262]=8'b01011111;
   assign rom_data[10263]=8'b01011011;
   assign rom_data[10264]=8'b01011110;
   assign rom_data[10265]=8'b01011001;
   assign rom_data[10266]=8'b01011110;
   assign rom_data[10267]=8'b01011000;
   assign rom_data[10268]=8'b01011110;
   assign rom_data[10269]=8'b01010111;
   assign rom_data[10270]=8'b01011110;
   assign rom_data[10271]=8'b01010101;
   assign rom_data[10272]=8'b01011110;
   assign rom_data[10273]=8'b01010100;
   assign rom_data[10274]=8'b01011110;
   assign rom_data[10275]=8'b01010010;
   assign rom_data[10276]=8'b01011110;
   assign rom_data[10277]=8'b01010001;
   assign rom_data[10278]=8'b01011110;
   assign rom_data[10279]=8'b01010000;
   assign rom_data[10280]=8'b01011110;
   assign rom_data[10281]=8'b01001110;
   assign rom_data[10282]=8'b01011110;
   assign rom_data[10283]=8'b01001101;
   assign rom_data[10284]=8'b01011110;
   assign rom_data[10285]=8'b01001100;
   assign rom_data[10286]=8'b01011110;
   assign rom_data[10287]=8'b01001010;
   assign rom_data[10288]=8'b01011110;
   assign rom_data[10289]=8'b01001001;
   assign rom_data[10290]=8'b01011110;
   assign rom_data[10291]=8'b01000111;
   assign rom_data[10292]=8'b01011110;
   assign rom_data[10293]=8'b01000110;
   assign rom_data[10294]=8'b01011110;
   assign rom_data[10295]=8'b01000101;
   assign rom_data[10296]=8'b01011110;
   assign rom_data[10297]=8'b01000100;
   assign rom_data[10298]=8'b01011110;
   assign rom_data[10299]=8'b01000010;
   assign rom_data[10300]=8'b01011110;
   assign rom_data[10301]=8'b01000001;
   assign rom_data[10302]=8'b01011110;
   assign rom_data[10303]=8'b01000000;
   assign rom_data[10304]=8'b01011110;
   assign rom_data[10305]=8'b00111110;
   assign rom_data[10306]=8'b01011110;
   assign rom_data[10307]=8'b00111101;
   assign rom_data[10308]=8'b01011110;
   assign rom_data[10309]=8'b00111100;
   assign rom_data[10310]=8'b01011110;
   assign rom_data[10311]=8'b00111011;
   assign rom_data[10312]=8'b01011110;
   assign rom_data[10313]=8'b00111010;
   assign rom_data[10314]=8'b01011110;
   assign rom_data[10315]=8'b00111001;
   assign rom_data[10316]=8'b01011110;
   assign rom_data[10317]=8'b00110111;
   assign rom_data[10318]=8'b01011110;
   assign rom_data[10319]=8'b00110110;
   assign rom_data[10320]=8'b01011110;
   assign rom_data[10321]=8'b00110101;
   assign rom_data[10322]=8'b01011110;
   assign rom_data[10323]=8'b00110100;
   assign rom_data[10324]=8'b01011110;
   assign rom_data[10325]=8'b00110011;
   assign rom_data[10326]=8'b01011110;
   assign rom_data[10327]=8'b00110011;
   assign rom_data[10328]=8'b01011110;
   assign rom_data[10329]=8'b00110010;
   assign rom_data[10330]=8'b01011110;
   assign rom_data[10331]=8'b00110001;
   assign rom_data[10332]=8'b01011110;
   assign rom_data[10333]=8'b00110000;
   assign rom_data[10334]=8'b01011110;
   assign rom_data[10335]=8'b00101111;
   assign rom_data[10336]=8'b01011110;
   assign rom_data[10337]=8'b00101111;
   assign rom_data[10338]=8'b01011110;
   assign rom_data[10339]=8'b00101110;
   assign rom_data[10340]=8'b01011101;
   assign rom_data[10341]=8'b00101110;
   assign rom_data[10342]=8'b01011101;
   assign rom_data[10343]=8'b00101101;
   assign rom_data[10344]=8'b01011101;
   assign rom_data[10345]=8'b00101101;
   assign rom_data[10346]=8'b01011101;
   assign rom_data[10347]=8'b00101100;
   assign rom_data[10348]=8'b01011101;
   assign rom_data[10349]=8'b00101100;
   assign rom_data[10350]=8'b01011101;
   assign rom_data[10351]=8'b00101100;
   assign rom_data[10352]=8'b01011101;
   assign rom_data[10353]=8'b00101100;
   assign rom_data[10354]=8'b01011101;
   assign rom_data[10355]=8'b00101100;
   assign rom_data[10356]=8'b01011101;
   assign rom_data[10357]=8'b00101100;
   assign rom_data[10358]=8'b01011101;
   assign rom_data[10359]=8'b00101100;
   assign rom_data[10360]=8'b01011101;
   assign rom_data[10361]=8'b00101101;
   assign rom_data[10362]=8'b01011101;
   assign rom_data[10363]=8'b00101101;
   assign rom_data[10364]=8'b01011101;
   assign rom_data[10365]=8'b00101101;
   assign rom_data[10366]=8'b01011101;
   assign rom_data[10367]=8'b00101110;
   assign rom_data[10368]=8'b01011101;
   assign rom_data[10369]=8'b00101111;
   assign rom_data[10370]=8'b01011101;
   assign rom_data[10371]=8'b00101111;
   assign rom_data[10372]=8'b01011101;
   assign rom_data[10373]=8'b00110000;
   assign rom_data[10374]=8'b01011101;
   assign rom_data[10375]=8'b00110001;
   assign rom_data[10376]=8'b01011101;
   assign rom_data[10377]=8'b00110001;
   assign rom_data[10378]=8'b01011101;
   assign rom_data[10379]=8'b00110010;
   assign rom_data[10380]=8'b01011101;
   assign rom_data[10381]=8'b00110011;
   assign rom_data[10382]=8'b01011101;
   assign rom_data[10383]=8'b00110100;
   assign rom_data[10384]=8'b01011101;
   assign rom_data[10385]=8'b00110101;
   assign rom_data[10386]=8'b01011101;
   assign rom_data[10387]=8'b00110110;
   assign rom_data[10388]=8'b01011101;
   assign rom_data[10389]=8'b00110111;
   assign rom_data[10390]=8'b01011101;
   assign rom_data[10391]=8'b00111000;
   assign rom_data[10392]=8'b01011101;
   assign rom_data[10393]=8'b00111010;
   assign rom_data[10394]=8'b01011101;
   assign rom_data[10395]=8'b00111011;
   assign rom_data[10396]=8'b01011101;
   assign rom_data[10397]=8'b00111100;
   assign rom_data[10398]=8'b01011101;
   assign rom_data[10399]=8'b00111101;
   assign rom_data[10400]=8'b01011101;
   assign rom_data[10401]=8'b00111110;
   assign rom_data[10402]=8'b01011101;
   assign rom_data[10403]=8'b01000000;
   assign rom_data[10404]=8'b01011101;
   assign rom_data[10405]=8'b01000001;
   assign rom_data[10406]=8'b01011101;
   assign rom_data[10407]=8'b01000010;
   assign rom_data[10408]=8'b01011100;
   assign rom_data[10409]=8'b01000100;
   assign rom_data[10410]=8'b01011100;
   assign rom_data[10411]=8'b01000101;
   assign rom_data[10412]=8'b01011100;
   assign rom_data[10413]=8'b01000110;
   assign rom_data[10414]=8'b01011100;
   assign rom_data[10415]=8'b01001000;
   assign rom_data[10416]=8'b01011100;
   assign rom_data[10417]=8'b01001001;
   assign rom_data[10418]=8'b01011100;
   assign rom_data[10419]=8'b01001010;
   assign rom_data[10420]=8'b01011100;
   assign rom_data[10421]=8'b01001100;
   assign rom_data[10422]=8'b01011100;
   assign rom_data[10423]=8'b01001101;
   assign rom_data[10424]=8'b01011100;
   assign rom_data[10425]=8'b01001110;
   assign rom_data[10426]=8'b01011100;
   assign rom_data[10427]=8'b01010000;
   assign rom_data[10428]=8'b01011100;
   assign rom_data[10429]=8'b01010001;
   assign rom_data[10430]=8'b01011100;
   assign rom_data[10431]=8'b01010011;
   assign rom_data[10432]=8'b01011100;
   assign rom_data[10433]=8'b01010100;
   assign rom_data[10434]=8'b01011100;
   assign rom_data[10435]=8'b01010101;
   assign rom_data[10436]=8'b01011100;
   assign rom_data[10437]=8'b01010111;
   assign rom_data[10438]=8'b01011100;
   assign rom_data[10439]=8'b01011000;
   assign rom_data[10440]=8'b01011100;
   assign rom_data[10441]=8'b01011010;
   assign rom_data[10442]=8'b01011100;
   assign rom_data[10443]=8'b01011011;
   assign rom_data[10444]=8'b01011100;
   assign rom_data[10445]=8'b01011100;
   assign rom_data[10446]=8'b01011100;
   assign rom_data[10447]=8'b01011110;
   assign rom_data[10448]=8'b01011100;
   assign rom_data[10449]=8'b01011111;
   assign rom_data[10450]=8'b01011100;
   assign rom_data[10451]=8'b01100001;
   assign rom_data[10452]=8'b01011100;
   assign rom_data[10453]=8'b01100010;
   assign rom_data[10454]=8'b01011100;
   assign rom_data[10455]=8'b01100011;
   assign rom_data[10456]=8'b01011100;
   assign rom_data[10457]=8'b01100101;
   assign rom_data[10458]=8'b01011100;
   assign rom_data[10459]=8'b01100110;
   assign rom_data[10460]=8'b01011100;
   assign rom_data[10461]=8'b01101000;
   assign rom_data[10462]=8'b01011100;
   assign rom_data[10463]=8'b01101001;
   assign rom_data[10464]=8'b01011100;
   assign rom_data[10465]=8'b01101010;
   assign rom_data[10466]=8'b01011100;
   assign rom_data[10467]=8'b01101100;
   assign rom_data[10468]=8'b01011100;
   assign rom_data[10469]=8'b01101101;
   assign rom_data[10470]=8'b01011100;
   assign rom_data[10471]=8'b01101110;
   assign rom_data[10472]=8'b01011100;
   assign rom_data[10473]=8'b01110000;
   assign rom_data[10474]=8'b01011100;
   assign rom_data[10475]=8'b01110001;
   assign rom_data[10476]=8'b01011100;
   assign rom_data[10477]=8'b01110010;
   assign rom_data[10478]=8'b01011100;
   assign rom_data[10479]=8'b01110100;
   assign rom_data[10480]=8'b01011100;
   assign rom_data[10481]=8'b01110101;
   assign rom_data[10482]=8'b01011100;
   assign rom_data[10483]=8'b01110110;
   assign rom_data[10484]=8'b01011100;
   assign rom_data[10485]=8'b01110111;
   assign rom_data[10486]=8'b01011100;
   assign rom_data[10487]=8'b01111001;
   assign rom_data[10488]=8'b01011100;
   assign rom_data[10489]=8'b01111010;
   assign rom_data[10490]=8'b01011100;
   assign rom_data[10491]=8'b01111011;
   assign rom_data[10492]=8'b01011011;
   assign rom_data[10493]=8'b01111100;
   assign rom_data[10494]=8'b01011011;
   assign rom_data[10495]=8'b01111101;
   assign rom_data[10496]=8'b01011011;
   assign rom_data[10497]=8'b01111110;
   assign rom_data[10498]=8'b01011011;
   assign rom_data[10499]=8'b01111111;
   assign rom_data[10500]=8'b01011011;
   assign rom_data[10501]=8'b10000000;
   assign rom_data[10502]=8'b01011011;
   assign rom_data[10503]=8'b10000001;
   assign rom_data[10504]=8'b01011011;
   assign rom_data[10505]=8'b10000010;
   assign rom_data[10506]=8'b01011011;
   assign rom_data[10507]=8'b10000011;
   assign rom_data[10508]=8'b01011011;
   assign rom_data[10509]=8'b10000100;
   assign rom_data[10510]=8'b01011011;
   assign rom_data[10511]=8'b10000101;
   assign rom_data[10512]=8'b01011011;
   assign rom_data[10513]=8'b10000110;
   assign rom_data[10514]=8'b01011011;
   assign rom_data[10515]=8'b10000110;
   assign rom_data[10516]=8'b01011011;
   assign rom_data[10517]=8'b10000111;
   assign rom_data[10518]=8'b01011011;
   assign rom_data[10519]=8'b10001000;
   assign rom_data[10520]=8'b01011011;
   assign rom_data[10521]=8'b10001000;
   assign rom_data[10522]=8'b01011011;
   assign rom_data[10523]=8'b10001001;
   assign rom_data[10524]=8'b01011011;
   assign rom_data[10525]=8'b10001001;
   assign rom_data[10526]=8'b01011011;
   assign rom_data[10527]=8'b10001001;
   assign rom_data[10528]=8'b01011011;
   assign rom_data[10529]=8'b10001010;
   assign rom_data[10530]=8'b01011011;
   assign rom_data[10531]=8'b10001010;
   assign rom_data[10532]=8'b01011011;
   assign rom_data[10533]=8'b10001010;
   assign rom_data[10534]=8'b01011011;
   assign rom_data[10535]=8'b10001010;
   assign rom_data[10536]=8'b01011011;
   assign rom_data[10537]=8'b10001010;
   assign rom_data[10538]=8'b01011011;
   assign rom_data[10539]=8'b10001001;
   assign rom_data[10540]=8'b01011011;
   assign rom_data[10541]=8'b10001001;
   assign rom_data[10542]=8'b01011011;
   assign rom_data[10543]=8'b10001001;
   assign rom_data[10544]=8'b01011011;
   assign rom_data[10545]=8'b10001000;
   assign rom_data[10546]=8'b01011011;
   assign rom_data[10547]=8'b10001000;
   assign rom_data[10548]=8'b01011011;
   assign rom_data[10549]=8'b10000111;
   assign rom_data[10550]=8'b01011011;
   assign rom_data[10551]=8'b10000111;
   assign rom_data[10552]=8'b01011011;
   assign rom_data[10553]=8'b10000110;
   assign rom_data[10554]=8'b01011011;
   assign rom_data[10555]=8'b10000101;
   assign rom_data[10556]=8'b01011011;
   assign rom_data[10557]=8'b10000100;
   assign rom_data[10558]=8'b01011010;
   assign rom_data[10559]=8'b10000011;
   assign rom_data[10560]=8'b01011010;
   assign rom_data[10561]=8'b10000011;
   assign rom_data[10562]=8'b01011010;
   assign rom_data[10563]=8'b10000010;
   assign rom_data[10564]=8'b01011010;
   assign rom_data[10565]=8'b10000001;
   assign rom_data[10566]=8'b01011010;
   assign rom_data[10567]=8'b10000000;
   assign rom_data[10568]=8'b01011010;
   assign rom_data[10569]=8'b01111110;
   assign rom_data[10570]=8'b01011010;
   assign rom_data[10571]=8'b01111101;
   assign rom_data[10572]=8'b01011010;
   assign rom_data[10573]=8'b01111100;
   assign rom_data[10574]=8'b01011010;
   assign rom_data[10575]=8'b01111011;
   assign rom_data[10576]=8'b01011010;
   assign rom_data[10577]=8'b01111010;
   assign rom_data[10578]=8'b01011010;
   assign rom_data[10579]=8'b01111001;
   assign rom_data[10580]=8'b01011010;
   assign rom_data[10581]=8'b01110111;
   assign rom_data[10582]=8'b01011010;
   assign rom_data[10583]=8'b01110110;
   assign rom_data[10584]=8'b01011010;
   assign rom_data[10585]=8'b01110101;
   assign rom_data[10586]=8'b01011010;
   assign rom_data[10587]=8'b01110100;
   assign rom_data[10588]=8'b01011010;
   assign rom_data[10589]=8'b01110010;
   assign rom_data[10590]=8'b01011010;
   assign rom_data[10591]=8'b01110001;
   assign rom_data[10592]=8'b01011010;
   assign rom_data[10593]=8'b01110000;
   assign rom_data[10594]=8'b01011010;
   assign rom_data[10595]=8'b01101110;
   assign rom_data[10596]=8'b01011010;
   assign rom_data[10597]=8'b01101101;
   assign rom_data[10598]=8'b01011010;
   assign rom_data[10599]=8'b01101100;
   assign rom_data[10600]=8'b01011010;
   assign rom_data[10601]=8'b01101010;
   assign rom_data[10602]=8'b01011010;
   assign rom_data[10603]=8'b01101001;
   assign rom_data[10604]=8'b01011010;
   assign rom_data[10605]=8'b01100111;
   assign rom_data[10606]=8'b01011010;
   assign rom_data[10607]=8'b01100110;
   assign rom_data[10608]=8'b01011010;
   assign rom_data[10609]=8'b01100101;
   assign rom_data[10610]=8'b01011010;
   assign rom_data[10611]=8'b01100011;
   assign rom_data[10612]=8'b01011010;
   assign rom_data[10613]=8'b01100010;
   assign rom_data[10614]=8'b01011010;
   assign rom_data[10615]=8'b01100000;
   assign rom_data[10616]=8'b01011010;
   assign rom_data[10617]=8'b01011111;
   assign rom_data[10618]=8'b01011010;
   assign rom_data[10619]=8'b01011110;
   assign rom_data[10620]=8'b01011010;
   assign rom_data[10621]=8'b01011100;
   assign rom_data[10622]=8'b01011010;
   assign rom_data[10623]=8'b01011011;
   assign rom_data[10624]=8'b01011010;
   assign rom_data[10625]=8'b01011001;
   assign rom_data[10626]=8'b01011010;
   assign rom_data[10627]=8'b01011000;
   assign rom_data[10628]=8'b01011010;
   assign rom_data[10629]=8'b01010111;
   assign rom_data[10630]=8'b01011010;
   assign rom_data[10631]=8'b01010101;
   assign rom_data[10632]=8'b01011010;
   assign rom_data[10633]=8'b01010100;
   assign rom_data[10634]=8'b01011010;
   assign rom_data[10635]=8'b01010010;
   assign rom_data[10636]=8'b01011010;
   assign rom_data[10637]=8'b01010001;
   assign rom_data[10638]=8'b01011010;
   assign rom_data[10639]=8'b01010000;
   assign rom_data[10640]=8'b01011001;
   assign rom_data[10641]=8'b01001110;
   assign rom_data[10642]=8'b01011001;
   assign rom_data[10643]=8'b01001101;
   assign rom_data[10644]=8'b01011001;
   assign rom_data[10645]=8'b01001100;
   assign rom_data[10646]=8'b01011001;
   assign rom_data[10647]=8'b01001010;
   assign rom_data[10648]=8'b01011001;
   assign rom_data[10649]=8'b01001001;
   assign rom_data[10650]=8'b01011001;
   assign rom_data[10651]=8'b01000111;
   assign rom_data[10652]=8'b01011001;
   assign rom_data[10653]=8'b01000110;
   assign rom_data[10654]=8'b01011001;
   assign rom_data[10655]=8'b01000101;
   assign rom_data[10656]=8'b01011001;
   assign rom_data[10657]=8'b01000100;
   assign rom_data[10658]=8'b01011001;
   assign rom_data[10659]=8'b01000010;
   assign rom_data[10660]=8'b01011001;
   assign rom_data[10661]=8'b01000001;
   assign rom_data[10662]=8'b01011001;
   assign rom_data[10663]=8'b01000000;
   assign rom_data[10664]=8'b01011001;
   assign rom_data[10665]=8'b00111110;
   assign rom_data[10666]=8'b01011001;
   assign rom_data[10667]=8'b00111101;
   assign rom_data[10668]=8'b01011001;
   assign rom_data[10669]=8'b00111100;
   assign rom_data[10670]=8'b01011001;
   assign rom_data[10671]=8'b00111011;
   assign rom_data[10672]=8'b01011001;
   assign rom_data[10673]=8'b00111010;
   assign rom_data[10674]=8'b01011001;
   assign rom_data[10675]=8'b00111001;
   assign rom_data[10676]=8'b01011001;
   assign rom_data[10677]=8'b00110111;
   assign rom_data[10678]=8'b01011001;
   assign rom_data[10679]=8'b00110110;
   assign rom_data[10680]=8'b01011001;
   assign rom_data[10681]=8'b00110101;
   assign rom_data[10682]=8'b01011001;
   assign rom_data[10683]=8'b00110100;
   assign rom_data[10684]=8'b01011001;
   assign rom_data[10685]=8'b00110011;
   assign rom_data[10686]=8'b01011001;
   assign rom_data[10687]=8'b00110011;
   assign rom_data[10688]=8'b01011001;
   assign rom_data[10689]=8'b00110010;
   assign rom_data[10690]=8'b01011001;
   assign rom_data[10691]=8'b00110001;
   assign rom_data[10692]=8'b01011001;
   assign rom_data[10693]=8'b00110000;
   assign rom_data[10694]=8'b01011001;
   assign rom_data[10695]=8'b00101111;
   assign rom_data[10696]=8'b01011001;
   assign rom_data[10697]=8'b00101111;
   assign rom_data[10698]=8'b01011001;
   assign rom_data[10699]=8'b00101110;
   assign rom_data[10700]=8'b01011001;
   assign rom_data[10701]=8'b00101110;
   assign rom_data[10702]=8'b01011001;
   assign rom_data[10703]=8'b00101101;
   assign rom_data[10704]=8'b01011001;
   assign rom_data[10705]=8'b00101101;
   assign rom_data[10706]=8'b01011001;
   assign rom_data[10707]=8'b00101100;
   assign rom_data[10708]=8'b01011001;
   assign rom_data[10709]=8'b00101100;
   assign rom_data[10710]=8'b01011001;
   assign rom_data[10711]=8'b00101100;
   assign rom_data[10712]=8'b01011000;
   assign rom_data[10713]=8'b00101100;
   assign rom_data[10714]=8'b01011000;
   assign rom_data[10715]=8'b00101100;
   assign rom_data[10716]=8'b01011000;
   assign rom_data[10717]=8'b00101100;
   assign rom_data[10718]=8'b01011000;
   assign rom_data[10719]=8'b00101100;
   assign rom_data[10720]=8'b01011000;
   assign rom_data[10721]=8'b00101101;
   assign rom_data[10722]=8'b01011000;
   assign rom_data[10723]=8'b00101101;
   assign rom_data[10724]=8'b01011000;
   assign rom_data[10725]=8'b00101101;
   assign rom_data[10726]=8'b01011000;
   assign rom_data[10727]=8'b00101110;
   assign rom_data[10728]=8'b01011000;
   assign rom_data[10729]=8'b00101111;
   assign rom_data[10730]=8'b01011000;
   assign rom_data[10731]=8'b00101111;
   assign rom_data[10732]=8'b01011000;
   assign rom_data[10733]=8'b00110000;
   assign rom_data[10734]=8'b01011000;
   assign rom_data[10735]=8'b00110001;
   assign rom_data[10736]=8'b01011000;
   assign rom_data[10737]=8'b00110001;
   assign rom_data[10738]=8'b01011000;
   assign rom_data[10739]=8'b00110010;
   assign rom_data[10740]=8'b01011000;
   assign rom_data[10741]=8'b00110011;
   assign rom_data[10742]=8'b01011000;
   assign rom_data[10743]=8'b00110100;
   assign rom_data[10744]=8'b01011000;
   assign rom_data[10745]=8'b00110101;
   assign rom_data[10746]=8'b01011000;
   assign rom_data[10747]=8'b00110110;
   assign rom_data[10748]=8'b01011000;
   assign rom_data[10749]=8'b00110111;
   assign rom_data[10750]=8'b01011000;
   assign rom_data[10751]=8'b00111000;
   assign rom_data[10752]=8'b01011000;
   assign rom_data[10753]=8'b00111010;
   assign rom_data[10754]=8'b01011000;
   assign rom_data[10755]=8'b00111011;
   assign rom_data[10756]=8'b01011000;
   assign rom_data[10757]=8'b00111100;
   assign rom_data[10758]=8'b01011000;
   assign rom_data[10759]=8'b00111101;
   assign rom_data[10760]=8'b01011000;
   assign rom_data[10761]=8'b00111110;
   assign rom_data[10762]=8'b01011000;
   assign rom_data[10763]=8'b01000000;
   assign rom_data[10764]=8'b01011000;
   assign rom_data[10765]=8'b01000001;
   assign rom_data[10766]=8'b01011000;
   assign rom_data[10767]=8'b01000010;
   assign rom_data[10768]=8'b01011000;
   assign rom_data[10769]=8'b01000100;
   assign rom_data[10770]=8'b01011000;
   assign rom_data[10771]=8'b01000101;
   assign rom_data[10772]=8'b01011000;
   assign rom_data[10773]=8'b01000110;
   assign rom_data[10774]=8'b01011000;
   assign rom_data[10775]=8'b01001000;
   assign rom_data[10776]=8'b01011000;
   assign rom_data[10777]=8'b01001001;
   assign rom_data[10778]=8'b01011000;
   assign rom_data[10779]=8'b01001010;
   assign rom_data[10780]=8'b01011000;
   assign rom_data[10781]=8'b01001100;
   assign rom_data[10782]=8'b01011000;
   assign rom_data[10783]=8'b01001101;
   assign rom_data[10784]=8'b01010111;
   assign rom_data[10785]=8'b01001110;
   assign rom_data[10786]=8'b01010111;
   assign rom_data[10787]=8'b01010000;
   assign rom_data[10788]=8'b01010111;
   assign rom_data[10789]=8'b01010001;
   assign rom_data[10790]=8'b01010111;
   assign rom_data[10791]=8'b01010011;
   assign rom_data[10792]=8'b01010111;
   assign rom_data[10793]=8'b01010100;
   assign rom_data[10794]=8'b01010111;
   assign rom_data[10795]=8'b01010101;
   assign rom_data[10796]=8'b01010111;
   assign rom_data[10797]=8'b01010111;
   assign rom_data[10798]=8'b01010111;
   assign rom_data[10799]=8'b01011000;
   assign rom_data[10800]=8'b01010111;
   assign rom_data[10801]=8'b01011010;
   assign rom_data[10802]=8'b01010111;
   assign rom_data[10803]=8'b01011011;
   assign rom_data[10804]=8'b01010111;
   assign rom_data[10805]=8'b01011100;
   assign rom_data[10806]=8'b01010111;
   assign rom_data[10807]=8'b01011110;
   assign rom_data[10808]=8'b01010111;
   assign rom_data[10809]=8'b01011111;
   assign rom_data[10810]=8'b01010111;
   assign rom_data[10811]=8'b01100001;
   assign rom_data[10812]=8'b01010111;
   assign rom_data[10813]=8'b01100010;
   assign rom_data[10814]=8'b01010111;
   assign rom_data[10815]=8'b01100011;
   assign rom_data[10816]=8'b01010111;
   assign rom_data[10817]=8'b01100101;
   assign rom_data[10818]=8'b01010111;
   assign rom_data[10819]=8'b01100110;
   assign rom_data[10820]=8'b01010111;
   assign rom_data[10821]=8'b01101000;
   assign rom_data[10822]=8'b01010111;
   assign rom_data[10823]=8'b01101001;
   assign rom_data[10824]=8'b01010111;
   assign rom_data[10825]=8'b01101010;
   assign rom_data[10826]=8'b01010111;
   assign rom_data[10827]=8'b01101100;
   assign rom_data[10828]=8'b01010111;
   assign rom_data[10829]=8'b01101101;
   assign rom_data[10830]=8'b01010111;
   assign rom_data[10831]=8'b01101110;
   assign rom_data[10832]=8'b01010111;
   assign rom_data[10833]=8'b01110000;
   assign rom_data[10834]=8'b01010111;
   assign rom_data[10835]=8'b01110001;
   assign rom_data[10836]=8'b01010111;
   assign rom_data[10837]=8'b01110010;
   assign rom_data[10838]=8'b01010111;
   assign rom_data[10839]=8'b01110100;
   assign rom_data[10840]=8'b01010111;
   assign rom_data[10841]=8'b01110101;
   assign rom_data[10842]=8'b01010111;
   assign rom_data[10843]=8'b01110110;
   assign rom_data[10844]=8'b01010111;
   assign rom_data[10845]=8'b01110111;
   assign rom_data[10846]=8'b01010111;
   assign rom_data[10847]=8'b01111001;
   assign rom_data[10848]=8'b01010111;
   assign rom_data[10849]=8'b01111010;
   assign rom_data[10850]=8'b01010111;
   assign rom_data[10851]=8'b01111011;
   assign rom_data[10852]=8'b01010111;
   assign rom_data[10853]=8'b01111100;
   assign rom_data[10854]=8'b01010111;
   assign rom_data[10855]=8'b01111101;
   assign rom_data[10856]=8'b01010111;
   assign rom_data[10857]=8'b01111110;
   assign rom_data[10858]=8'b01010111;
   assign rom_data[10859]=8'b01111111;
   assign rom_data[10860]=8'b01010111;
   assign rom_data[10861]=8'b10000000;
   assign rom_data[10862]=8'b01010111;
   assign rom_data[10863]=8'b10000001;
   assign rom_data[10864]=8'b01010111;
   assign rom_data[10865]=8'b10000010;
   assign rom_data[10866]=8'b01010110;
   assign rom_data[10867]=8'b10000011;
   assign rom_data[10868]=8'b01010110;
   assign rom_data[10869]=8'b10000100;
   assign rom_data[10870]=8'b01010110;
   assign rom_data[10871]=8'b10000101;
   assign rom_data[10872]=8'b01010110;
   assign rom_data[10873]=8'b10000110;
   assign rom_data[10874]=8'b01010110;
   assign rom_data[10875]=8'b10000110;
   assign rom_data[10876]=8'b01010110;
   assign rom_data[10877]=8'b10000111;
   assign rom_data[10878]=8'b01010110;
   assign rom_data[10879]=8'b10001000;
   assign rom_data[10880]=8'b01010110;
   assign rom_data[10881]=8'b10001000;
   assign rom_data[10882]=8'b01010110;
   assign rom_data[10883]=8'b10001001;
   assign rom_data[10884]=8'b01010110;
   assign rom_data[10885]=8'b10001001;
   assign rom_data[10886]=8'b01010110;
   assign rom_data[10887]=8'b10001001;
   assign rom_data[10888]=8'b01010110;
   assign rom_data[10889]=8'b10001010;
   assign rom_data[10890]=8'b01010110;
   assign rom_data[10891]=8'b10001010;
   assign rom_data[10892]=8'b01010110;
   assign rom_data[10893]=8'b10001010;
   assign rom_data[10894]=8'b01010110;
   assign rom_data[10895]=8'b10001010;
   assign rom_data[10896]=8'b01010110;
   assign rom_data[10897]=8'b10001010;
   assign rom_data[10898]=8'b01010110;
   assign rom_data[10899]=8'b10001001;
   assign rom_data[10900]=8'b01010110;
   assign rom_data[10901]=8'b10001001;
   assign rom_data[10902]=8'b01010110;
   assign rom_data[10903]=8'b10001001;
   assign rom_data[10904]=8'b01010110;
   assign rom_data[10905]=8'b10001000;
   assign rom_data[10906]=8'b01010110;
   assign rom_data[10907]=8'b10001000;
   assign rom_data[10908]=8'b01010110;
   assign rom_data[10909]=8'b10000111;
   assign rom_data[10910]=8'b01010110;
   assign rom_data[10911]=8'b10000111;
   assign rom_data[10912]=8'b01010110;
   assign rom_data[10913]=8'b10000110;
   assign rom_data[10914]=8'b01010110;
   assign rom_data[10915]=8'b10000101;
   assign rom_data[10916]=8'b01010110;
   assign rom_data[10917]=8'b10000100;
   assign rom_data[10918]=8'b01010110;
   assign rom_data[10919]=8'b10000011;
   assign rom_data[10920]=8'b01010110;
   assign rom_data[10921]=8'b10000011;
   assign rom_data[10922]=8'b01010110;
   assign rom_data[10923]=8'b10000010;
   assign rom_data[10924]=8'b01010110;
   assign rom_data[10925]=8'b10000001;
   assign rom_data[10926]=8'b01010110;
   assign rom_data[10927]=8'b10000000;
   assign rom_data[10928]=8'b01010110;
   assign rom_data[10929]=8'b01111110;
   assign rom_data[10930]=8'b01010110;
   assign rom_data[10931]=8'b01111101;
   assign rom_data[10932]=8'b01010101;
   assign rom_data[10933]=8'b01111100;
   assign rom_data[10934]=8'b01010101;
   assign rom_data[10935]=8'b01111011;
   assign rom_data[10936]=8'b01010101;
   assign rom_data[10937]=8'b01111010;
   assign rom_data[10938]=8'b01010101;
   assign rom_data[10939]=8'b01111001;
   assign rom_data[10940]=8'b01010101;
   assign rom_data[10941]=8'b01110111;
   assign rom_data[10942]=8'b01010101;
   assign rom_data[10943]=8'b01110110;
   assign rom_data[10944]=8'b01010101;
   assign rom_data[10945]=8'b01110101;
   assign rom_data[10946]=8'b01010101;
   assign rom_data[10947]=8'b01110100;
   assign rom_data[10948]=8'b01010101;
   assign rom_data[10949]=8'b01110010;
   assign rom_data[10950]=8'b01010101;
   assign rom_data[10951]=8'b01110001;
   assign rom_data[10952]=8'b01010101;
   assign rom_data[10953]=8'b01110000;
   assign rom_data[10954]=8'b01010101;
   assign rom_data[10955]=8'b01101110;
   assign rom_data[10956]=8'b01010101;
   assign rom_data[10957]=8'b01101101;
   assign rom_data[10958]=8'b01010101;
   assign rom_data[10959]=8'b01101100;
   assign rom_data[10960]=8'b01010101;
   assign rom_data[10961]=8'b01101010;
   assign rom_data[10962]=8'b01010101;
   assign rom_data[10963]=8'b01101001;
   assign rom_data[10964]=8'b01010101;
   assign rom_data[10965]=8'b01100111;
   assign rom_data[10966]=8'b01010101;
   assign rom_data[10967]=8'b01100110;
   assign rom_data[10968]=8'b01010101;
   assign rom_data[10969]=8'b01100101;
   assign rom_data[10970]=8'b01010101;
   assign rom_data[10971]=8'b01100011;
   assign rom_data[10972]=8'b01010101;
   assign rom_data[10973]=8'b01100010;
   assign rom_data[10974]=8'b01010101;
   assign rom_data[10975]=8'b01100000;
   assign rom_data[10976]=8'b01010101;
   assign rom_data[10977]=8'b01011111;
   assign rom_data[10978]=8'b01010101;
   assign rom_data[10979]=8'b01011110;
   assign rom_data[10980]=8'b01010101;
   assign rom_data[10981]=8'b01011100;
   assign rom_data[10982]=8'b01010101;
   assign rom_data[10983]=8'b01011011;
   assign rom_data[10984]=8'b01010101;
   assign rom_data[10985]=8'b01011001;
   assign rom_data[10986]=8'b01010101;
   assign rom_data[10987]=8'b01011000;
   assign rom_data[10988]=8'b01010101;
   assign rom_data[10989]=8'b01010111;
   assign rom_data[10990]=8'b01010101;
   assign rom_data[10991]=8'b01010101;
   assign rom_data[10992]=8'b01010101;
   assign rom_data[10993]=8'b01010100;
   assign rom_data[10994]=8'b01010101;
   assign rom_data[10995]=8'b01010010;
   assign rom_data[10996]=8'b01010101;
   assign rom_data[10997]=8'b01010001;
   assign rom_data[10998]=8'b01010101;
   assign rom_data[10999]=8'b01010000;
   assign rom_data[11000]=8'b01010101;
   assign rom_data[11001]=8'b01001110;
   assign rom_data[11002]=8'b01010101;
   assign rom_data[11003]=8'b01001101;
   assign rom_data[11004]=8'b01010101;
   assign rom_data[11005]=8'b01001100;
   assign rom_data[11006]=8'b01010101;
   assign rom_data[11007]=8'b01001010;
   assign rom_data[11008]=8'b01010101;
   assign rom_data[11009]=8'b01001001;
   assign rom_data[11010]=8'b01010101;
   assign rom_data[11011]=8'b01000111;
   assign rom_data[11012]=8'b01010101;
   assign rom_data[11013]=8'b01000110;
   assign rom_data[11014]=8'b01010101;
   assign rom_data[11015]=8'b01000101;
   assign rom_data[11016]=8'b01010100;
   assign rom_data[11017]=8'b01000100;
   assign rom_data[11018]=8'b01010100;
   assign rom_data[11019]=8'b01000010;
   assign rom_data[11020]=8'b01010100;
   assign rom_data[11021]=8'b01000001;
   assign rom_data[11022]=8'b01010100;
   assign rom_data[11023]=8'b01000000;
   assign rom_data[11024]=8'b01010100;
   assign rom_data[11025]=8'b00111110;
   assign rom_data[11026]=8'b01010100;
   assign rom_data[11027]=8'b00111101;
   assign rom_data[11028]=8'b01010100;
   assign rom_data[11029]=8'b00111100;
   assign rom_data[11030]=8'b01010100;
   assign rom_data[11031]=8'b00111011;
   assign rom_data[11032]=8'b01010100;
   assign rom_data[11033]=8'b00111010;
   assign rom_data[11034]=8'b01010100;
   assign rom_data[11035]=8'b00111001;
   assign rom_data[11036]=8'b01010100;
   assign rom_data[11037]=8'b00110111;
   assign rom_data[11038]=8'b01010100;
   assign rom_data[11039]=8'b00110110;
   assign rom_data[11040]=8'b01010100;
   assign rom_data[11041]=8'b00110101;
   assign rom_data[11042]=8'b01010100;
   assign rom_data[11043]=8'b00110100;
   assign rom_data[11044]=8'b01010100;
   assign rom_data[11045]=8'b00110011;
   assign rom_data[11046]=8'b01010100;
   assign rom_data[11047]=8'b00110011;
   assign rom_data[11048]=8'b01010100;
   assign rom_data[11049]=8'b00110010;
   assign rom_data[11050]=8'b01010100;
   assign rom_data[11051]=8'b00110001;
   assign rom_data[11052]=8'b01010100;
   assign rom_data[11053]=8'b00110000;
   assign rom_data[11054]=8'b01010100;
   assign rom_data[11055]=8'b00101111;
   assign rom_data[11056]=8'b01010100;
   assign rom_data[11057]=8'b00101111;
   assign rom_data[11058]=8'b01010100;
   assign rom_data[11059]=8'b00101110;
   assign rom_data[11060]=8'b01010100;
   assign rom_data[11061]=8'b00101110;
   assign rom_data[11062]=8'b01010100;
   assign rom_data[11063]=8'b00101101;
   assign rom_data[11064]=8'b01010100;
   assign rom_data[11065]=8'b00101101;
   assign rom_data[11066]=8'b01010100;
   assign rom_data[11067]=8'b00101100;
   assign rom_data[11068]=8'b01010100;
   assign rom_data[11069]=8'b00101100;
   assign rom_data[11070]=8'b01010100;
   assign rom_data[11071]=8'b00101100;
   assign rom_data[11072]=8'b01010100;
   assign rom_data[11073]=8'b00101100;
   assign rom_data[11074]=8'b01010100;
   assign rom_data[11075]=8'b00101100;
   assign rom_data[11076]=8'b01010100;
   assign rom_data[11077]=8'b00101100;
   assign rom_data[11078]=8'b01010100;
   assign rom_data[11079]=8'b00101100;
   assign rom_data[11080]=8'b01010100;
   assign rom_data[11081]=8'b00101101;
   assign rom_data[11082]=8'b01010100;
   assign rom_data[11083]=8'b00101101;
   assign rom_data[11084]=8'b01010011;
   assign rom_data[11085]=8'b00101101;
   assign rom_data[11086]=8'b01010011;
   assign rom_data[11087]=8'b00101110;
   assign rom_data[11088]=8'b01010011;
   assign rom_data[11089]=8'b00101111;
   assign rom_data[11090]=8'b01010011;
   assign rom_data[11091]=8'b00101111;
   assign rom_data[11092]=8'b01010011;
   assign rom_data[11093]=8'b00110000;
   assign rom_data[11094]=8'b01010011;
   assign rom_data[11095]=8'b00110001;
   assign rom_data[11096]=8'b01010011;
   assign rom_data[11097]=8'b00110010;
   assign rom_data[11098]=8'b01010011;
   assign rom_data[11099]=8'b00110010;
   assign rom_data[11100]=8'b01010011;
   assign rom_data[11101]=8'b00110011;
   assign rom_data[11102]=8'b01010011;
   assign rom_data[11103]=8'b00110100;
   assign rom_data[11104]=8'b01010011;
   assign rom_data[11105]=8'b00110101;
   assign rom_data[11106]=8'b01010011;
   assign rom_data[11107]=8'b00110110;
   assign rom_data[11108]=8'b01010011;
   assign rom_data[11109]=8'b00110111;
   assign rom_data[11110]=8'b01010011;
   assign rom_data[11111]=8'b00111001;
   assign rom_data[11112]=8'b01010011;
   assign rom_data[11113]=8'b00111010;
   assign rom_data[11114]=8'b01010011;
   assign rom_data[11115]=8'b00111011;
   assign rom_data[11116]=8'b01010011;
   assign rom_data[11117]=8'b00111100;
   assign rom_data[11118]=8'b01010011;
   assign rom_data[11119]=8'b00111101;
   assign rom_data[11120]=8'b01010011;
   assign rom_data[11121]=8'b00111110;
   assign rom_data[11122]=8'b01010011;
   assign rom_data[11123]=8'b01000000;
   assign rom_data[11124]=8'b01010011;
   assign rom_data[11125]=8'b01000001;
   assign rom_data[11126]=8'b01010011;
   assign rom_data[11127]=8'b01000010;
   assign rom_data[11128]=8'b01010011;
   assign rom_data[11129]=8'b01000100;
   assign rom_data[11130]=8'b01010011;
   assign rom_data[11131]=8'b01000101;
   assign rom_data[11132]=8'b01010011;
   assign rom_data[11133]=8'b01000110;
   assign rom_data[11134]=8'b01010011;
   assign rom_data[11135]=8'b01001000;
   assign rom_data[11136]=8'b01010011;
   assign rom_data[11137]=8'b01001001;
   assign rom_data[11138]=8'b01010011;
   assign rom_data[11139]=8'b01001010;
   assign rom_data[11140]=8'b01010011;
   assign rom_data[11141]=8'b01001100;
   assign rom_data[11142]=8'b01010011;
   assign rom_data[11143]=8'b01001101;
   assign rom_data[11144]=8'b01010011;
   assign rom_data[11145]=8'b01001110;
   assign rom_data[11146]=8'b01010011;
   assign rom_data[11147]=8'b01010000;
   assign rom_data[11148]=8'b01010011;
   assign rom_data[11149]=8'b01010001;
   assign rom_data[11150]=8'b01010011;
   assign rom_data[11151]=8'b01010011;
   assign rom_data[11152]=8'b01010011;
   assign rom_data[11153]=8'b01010100;
   assign rom_data[11154]=8'b01010011;
   assign rom_data[11155]=8'b01010101;
   assign rom_data[11156]=8'b01010011;
   assign rom_data[11157]=8'b01010111;
   assign rom_data[11158]=8'b01010011;
   assign rom_data[11159]=8'b01011000;
   assign rom_data[11160]=8'b01010011;
   assign rom_data[11161]=8'b01011010;
   assign rom_data[11162]=8'b01010010;
   assign rom_data[11163]=8'b01011011;
   assign rom_data[11164]=8'b01010010;
   assign rom_data[11165]=8'b01011100;
   assign rom_data[11166]=8'b01010010;
   assign rom_data[11167]=8'b01011110;
   assign rom_data[11168]=8'b01010010;
   assign rom_data[11169]=8'b01011111;
   assign rom_data[11170]=8'b01010010;
   assign rom_data[11171]=8'b01100001;
   assign rom_data[11172]=8'b01010010;
   assign rom_data[11173]=8'b01100010;
   assign rom_data[11174]=8'b01010010;
   assign rom_data[11175]=8'b01100011;
   assign rom_data[11176]=8'b01010010;
   assign rom_data[11177]=8'b01100101;
   assign rom_data[11178]=8'b01010010;
   assign rom_data[11179]=8'b01100110;
   assign rom_data[11180]=8'b01010010;
   assign rom_data[11181]=8'b01101000;
   assign rom_data[11182]=8'b01010010;
   assign rom_data[11183]=8'b01101001;
   assign rom_data[11184]=8'b01010010;
   assign rom_data[11185]=8'b01101010;
   assign rom_data[11186]=8'b01010010;
   assign rom_data[11187]=8'b01101100;
   assign rom_data[11188]=8'b01010010;
   assign rom_data[11189]=8'b01101101;
   assign rom_data[11190]=8'b01010010;
   assign rom_data[11191]=8'b01101110;
   assign rom_data[11192]=8'b01010010;
   assign rom_data[11193]=8'b01110000;
   assign rom_data[11194]=8'b01010010;
   assign rom_data[11195]=8'b01110001;
   assign rom_data[11196]=8'b01010010;
   assign rom_data[11197]=8'b01110010;
   assign rom_data[11198]=8'b01010010;
   assign rom_data[11199]=8'b01110100;
   assign rom_data[11200]=8'b01010010;
   assign rom_data[11201]=8'b01110101;
   assign rom_data[11202]=8'b01010010;
   assign rom_data[11203]=8'b01110110;
   assign rom_data[11204]=8'b01010010;
   assign rom_data[11205]=8'b01110111;
   assign rom_data[11206]=8'b01010010;
   assign rom_data[11207]=8'b01111001;
   assign rom_data[11208]=8'b01010010;
   assign rom_data[11209]=8'b01111010;
   assign rom_data[11210]=8'b01010010;
   assign rom_data[11211]=8'b01111011;
   assign rom_data[11212]=8'b01010010;
   assign rom_data[11213]=8'b01111100;
   assign rom_data[11214]=8'b01010010;
   assign rom_data[11215]=8'b01111101;
   assign rom_data[11216]=8'b01010010;
   assign rom_data[11217]=8'b01111110;
   assign rom_data[11218]=8'b01010010;
   assign rom_data[11219]=8'b01111111;
   assign rom_data[11220]=8'b01010010;
   assign rom_data[11221]=8'b10000000;
   assign rom_data[11222]=8'b01010010;
   assign rom_data[11223]=8'b10000001;
   assign rom_data[11224]=8'b01010010;
   assign rom_data[11225]=8'b10000010;
   assign rom_data[11226]=8'b01010010;
   assign rom_data[11227]=8'b10000011;
   assign rom_data[11228]=8'b01010010;
   assign rom_data[11229]=8'b10000100;
   assign rom_data[11230]=8'b01010010;
   assign rom_data[11231]=8'b10000101;
   assign rom_data[11232]=8'b01010010;
   assign rom_data[11233]=8'b10000110;
   assign rom_data[11234]=8'b01010010;
   assign rom_data[11235]=8'b10000110;
   assign rom_data[11236]=8'b01010010;
   assign rom_data[11237]=8'b10000111;
   assign rom_data[11238]=8'b01010001;
   assign rom_data[11239]=8'b10001000;
   assign rom_data[11240]=8'b01010001;
   assign rom_data[11241]=8'b10001000;
   assign rom_data[11242]=8'b01010001;
   assign rom_data[11243]=8'b10001001;
   assign rom_data[11244]=8'b01010001;
   assign rom_data[11245]=8'b10001001;
   assign rom_data[11246]=8'b01010001;
   assign rom_data[11247]=8'b10001001;
   assign rom_data[11248]=8'b01010001;
   assign rom_data[11249]=8'b10001010;
   assign rom_data[11250]=8'b01010001;
   assign rom_data[11251]=8'b10001010;
   assign rom_data[11252]=8'b01010001;
   assign rom_data[11253]=8'b10001010;
   assign rom_data[11254]=8'b01010001;
   assign rom_data[11255]=8'b10001010;
   assign rom_data[11256]=8'b01010001;
   assign rom_data[11257]=8'b10001010;
   assign rom_data[11258]=8'b01010001;
   assign rom_data[11259]=8'b10001001;
   assign rom_data[11260]=8'b01010001;
   assign rom_data[11261]=8'b10001001;
   assign rom_data[11262]=8'b01010001;
   assign rom_data[11263]=8'b10001001;
   assign rom_data[11264]=8'b01010001;
   assign rom_data[11265]=8'b10001000;
   assign rom_data[11266]=8'b01010001;
   assign rom_data[11267]=8'b10001000;
   assign rom_data[11268]=8'b01010001;
   assign rom_data[11269]=8'b10000111;
   assign rom_data[11270]=8'b01010001;
   assign rom_data[11271]=8'b10000111;
   assign rom_data[11272]=8'b01010001;
   assign rom_data[11273]=8'b10000110;
   assign rom_data[11274]=8'b01010001;
   assign rom_data[11275]=8'b10000101;
   assign rom_data[11276]=8'b01010001;
   assign rom_data[11277]=8'b10000100;
   assign rom_data[11278]=8'b01010001;
   assign rom_data[11279]=8'b10000011;
   assign rom_data[11280]=8'b01010001;
   assign rom_data[11281]=8'b10000011;
   assign rom_data[11282]=8'b01010001;
   assign rom_data[11283]=8'b10000010;
   assign rom_data[11284]=8'b01010001;
   assign rom_data[11285]=8'b10000001;
   assign rom_data[11286]=8'b01010001;
   assign rom_data[11287]=8'b10000000;
   assign rom_data[11288]=8'b01010001;
   assign rom_data[11289]=8'b01111110;
   assign rom_data[11290]=8'b01010001;
   assign rom_data[11291]=8'b01111101;
   assign rom_data[11292]=8'b01010001;
   assign rom_data[11293]=8'b01111100;
   assign rom_data[11294]=8'b01010001;
   assign rom_data[11295]=8'b01111011;
   assign rom_data[11296]=8'b01010001;
   assign rom_data[11297]=8'b01111010;
   assign rom_data[11298]=8'b01010001;
   assign rom_data[11299]=8'b01111001;
   assign rom_data[11300]=8'b01010001;
   assign rom_data[11301]=8'b01110111;
   assign rom_data[11302]=8'b01010001;
   assign rom_data[11303]=8'b01110110;
   assign rom_data[11304]=8'b01010001;
   assign rom_data[11305]=8'b01110101;
   assign rom_data[11306]=8'b01010000;
   assign rom_data[11307]=8'b01110100;
   assign rom_data[11308]=8'b01010000;
   assign rom_data[11309]=8'b01110010;
   assign rom_data[11310]=8'b01010000;
   assign rom_data[11311]=8'b01110001;
   assign rom_data[11312]=8'b01010000;
   assign rom_data[11313]=8'b01110000;
   assign rom_data[11314]=8'b01010000;
   assign rom_data[11315]=8'b01101110;
   assign rom_data[11316]=8'b01010000;
   assign rom_data[11317]=8'b01101101;
   assign rom_data[11318]=8'b01010000;
   assign rom_data[11319]=8'b01101100;
   assign rom_data[11320]=8'b01010000;
   assign rom_data[11321]=8'b01101010;
   assign rom_data[11322]=8'b01010000;
   assign rom_data[11323]=8'b01101001;
   assign rom_data[11324]=8'b01010000;
   assign rom_data[11325]=8'b01100111;
   assign rom_data[11326]=8'b01010000;
   assign rom_data[11327]=8'b01100110;
   assign rom_data[11328]=8'b01010000;
   assign rom_data[11329]=8'b01100101;
   assign rom_data[11330]=8'b01010000;
   assign rom_data[11331]=8'b01100011;
   assign rom_data[11332]=8'b01010000;
   assign rom_data[11333]=8'b01100010;
   assign rom_data[11334]=8'b01010000;
   assign rom_data[11335]=8'b01100000;
   assign rom_data[11336]=8'b01010000;
   assign rom_data[11337]=8'b01011111;
   assign rom_data[11338]=8'b01010000;
   assign rom_data[11339]=8'b01011110;
   assign rom_data[11340]=8'b01010000;
   assign rom_data[11341]=8'b01011100;
   assign rom_data[11342]=8'b01010000;
   assign rom_data[11343]=8'b01011011;
   assign rom_data[11344]=8'b01010000;
   assign rom_data[11345]=8'b01011001;
   assign rom_data[11346]=8'b01010000;
   assign rom_data[11347]=8'b01011000;
   assign rom_data[11348]=8'b01010000;
   assign rom_data[11349]=8'b01010111;
   assign rom_data[11350]=8'b01010000;
   assign rom_data[11351]=8'b01010101;
   assign rom_data[11352]=8'b01010000;
   assign rom_data[11353]=8'b01010100;
   assign rom_data[11354]=8'b01010000;
   assign rom_data[11355]=8'b01010010;
   assign rom_data[11356]=8'b01010000;
   assign rom_data[11357]=8'b01010001;
   assign rom_data[11358]=8'b01010000;
   assign rom_data[11359]=8'b01010000;
   assign rom_data[11360]=8'b01010000;
   assign rom_data[11361]=8'b01001110;
   assign rom_data[11362]=8'b01010000;
   assign rom_data[11363]=8'b01001101;
   assign rom_data[11364]=8'b01010000;
   assign rom_data[11365]=8'b01001100;
   assign rom_data[11366]=8'b01010000;
   assign rom_data[11367]=8'b01001010;
   assign rom_data[11368]=8'b01010000;
   assign rom_data[11369]=8'b01001001;
   assign rom_data[11370]=8'b01010000;
   assign rom_data[11371]=8'b01000111;
   assign rom_data[11372]=8'b01010000;
   assign rom_data[11373]=8'b01000110;
   assign rom_data[11374]=8'b01010000;
   assign rom_data[11375]=8'b01000101;
   assign rom_data[11376]=8'b01010000;
   assign rom_data[11377]=8'b01000100;
   assign rom_data[11378]=8'b01010000;
   assign rom_data[11379]=8'b01000010;
   assign rom_data[11380]=8'b01010000;
   assign rom_data[11381]=8'b01000001;
   assign rom_data[11382]=8'b01010000;
   assign rom_data[11383]=8'b01000000;
   assign rom_data[11384]=8'b01010000;
   assign rom_data[11385]=8'b00111110;
   assign rom_data[11386]=8'b01010000;
   assign rom_data[11387]=8'b00111101;
   assign rom_data[11388]=8'b01010000;
   assign rom_data[11389]=8'b00111100;
   assign rom_data[11390]=8'b01001111;
   assign rom_data[11391]=8'b00111011;
   assign rom_data[11392]=8'b01001111;
   assign rom_data[11393]=8'b00111010;
   assign rom_data[11394]=8'b01001111;
   assign rom_data[11395]=8'b00111001;
   assign rom_data[11396]=8'b01001111;
   assign rom_data[11397]=8'b00110111;
   assign rom_data[11398]=8'b01001111;
   assign rom_data[11399]=8'b00110110;
   assign rom_data[11400]=8'b01001111;
   assign rom_data[11401]=8'b00110101;
   assign rom_data[11402]=8'b01001111;
   assign rom_data[11403]=8'b00110100;
   assign rom_data[11404]=8'b01001111;
   assign rom_data[11405]=8'b00110011;
   assign rom_data[11406]=8'b01001111;
   assign rom_data[11407]=8'b00110011;
   assign rom_data[11408]=8'b01001111;
   assign rom_data[11409]=8'b00110010;
   assign rom_data[11410]=8'b01001111;
   assign rom_data[11411]=8'b00110001;
   assign rom_data[11412]=8'b01001111;
   assign rom_data[11413]=8'b00110000;
   assign rom_data[11414]=8'b01001111;
   assign rom_data[11415]=8'b00101111;
   assign rom_data[11416]=8'b01001111;
   assign rom_data[11417]=8'b00101111;
   assign rom_data[11418]=8'b01001111;
   assign rom_data[11419]=8'b00101110;
   assign rom_data[11420]=8'b01001111;
   assign rom_data[11421]=8'b00101110;
   assign rom_data[11422]=8'b01001111;
   assign rom_data[11423]=8'b00101101;
   assign rom_data[11424]=8'b01001111;
   assign rom_data[11425]=8'b00101101;
   assign rom_data[11426]=8'b01001111;
   assign rom_data[11427]=8'b00101100;
   assign rom_data[11428]=8'b01001111;
   assign rom_data[11429]=8'b00101100;
   assign rom_data[11430]=8'b01001111;
   assign rom_data[11431]=8'b00101100;
   assign rom_data[11432]=8'b01001111;
   assign rom_data[11433]=8'b00101100;
   assign rom_data[11434]=8'b01001111;
   assign rom_data[11435]=8'b00101100;
   assign rom_data[11436]=8'b01001111;
   assign rom_data[11437]=8'b00101100;
   assign rom_data[11438]=8'b01001111;
   assign rom_data[11439]=8'b00101100;
   assign rom_data[11440]=8'b01001111;
   assign rom_data[11441]=8'b00101101;
   assign rom_data[11442]=8'b01001111;
   assign rom_data[11443]=8'b00101101;
   assign rom_data[11444]=8'b01001111;
   assign rom_data[11445]=8'b00101101;
   assign rom_data[11446]=8'b01001111;
   assign rom_data[11447]=8'b00101110;
   assign rom_data[11448]=8'b01001111;
   assign rom_data[11449]=8'b00101111;
   assign rom_data[11450]=8'b01001111;
   assign rom_data[11451]=8'b00101111;
   assign rom_data[11452]=8'b01001111;
   assign rom_data[11453]=8'b00110000;
   assign rom_data[11454]=8'b01001111;
   assign rom_data[11455]=8'b00110001;
   assign rom_data[11456]=8'b01001110;
   assign rom_data[11457]=8'b00110010;
   assign rom_data[11458]=8'b01001110;
   assign rom_data[11459]=8'b00110010;
   assign rom_data[11460]=8'b01001110;
   assign rom_data[11461]=8'b00110011;
   assign rom_data[11462]=8'b01001110;
   assign rom_data[11463]=8'b00110100;
   assign rom_data[11464]=8'b01001110;
   assign rom_data[11465]=8'b00110101;
   assign rom_data[11466]=8'b01001110;
   assign rom_data[11467]=8'b00110110;
   assign rom_data[11468]=8'b01001110;
   assign rom_data[11469]=8'b00110111;
   assign rom_data[11470]=8'b01001110;
   assign rom_data[11471]=8'b00111001;
   assign rom_data[11472]=8'b01001110;
   assign rom_data[11473]=8'b00111010;
   assign rom_data[11474]=8'b01001110;
   assign rom_data[11475]=8'b00111011;
   assign rom_data[11476]=8'b01001110;
   assign rom_data[11477]=8'b00111100;
   assign rom_data[11478]=8'b01001110;
   assign rom_data[11479]=8'b00111101;
   assign rom_data[11480]=8'b01001110;
   assign rom_data[11481]=8'b00111110;
   assign rom_data[11482]=8'b01001110;
   assign rom_data[11483]=8'b01000000;
   assign rom_data[11484]=8'b01001110;
   assign rom_data[11485]=8'b01000001;
   assign rom_data[11486]=8'b01001110;
   assign rom_data[11487]=8'b01000010;
   assign rom_data[11488]=8'b01001110;
   assign rom_data[11489]=8'b01000100;
   assign rom_data[11490]=8'b01001110;
   assign rom_data[11491]=8'b01000101;
   assign rom_data[11492]=8'b01001110;
   assign rom_data[11493]=8'b01000110;
   assign rom_data[11494]=8'b01001110;
   assign rom_data[11495]=8'b01001000;
   assign rom_data[11496]=8'b01001110;
   assign rom_data[11497]=8'b01001001;
   assign rom_data[11498]=8'b01001110;
   assign rom_data[11499]=8'b01001010;
   assign rom_data[11500]=8'b01001110;
   assign rom_data[11501]=8'b01001100;
   assign rom_data[11502]=8'b01001110;
   assign rom_data[11503]=8'b01001101;
   assign rom_data[11504]=8'b01001110;
   assign rom_data[11505]=8'b01001110;
   assign rom_data[11506]=8'b01001110;
   assign rom_data[11507]=8'b01010000;
   assign rom_data[11508]=8'b01001110;
   assign rom_data[11509]=8'b01010001;
   assign rom_data[11510]=8'b01001110;
   assign rom_data[11511]=8'b01010011;
   assign rom_data[11512]=8'b01001110;
   assign rom_data[11513]=8'b01010100;
   assign rom_data[11514]=8'b01001110;
   assign rom_data[11515]=8'b01010101;
   assign rom_data[11516]=8'b01001110;
   assign rom_data[11517]=8'b01010111;
   assign rom_data[11518]=8'b01001110;
   assign rom_data[11519]=8'b01011000;
   assign rom_data[11520]=8'b01001110;
   assign rom_data[11521]=8'b01011010;
   assign rom_data[11522]=8'b01001110;
   assign rom_data[11523]=8'b01011011;
   assign rom_data[11524]=8'b01001110;
   assign rom_data[11525]=8'b01011100;
   assign rom_data[11526]=8'b01001110;
   assign rom_data[11527]=8'b01011110;
   assign rom_data[11528]=8'b01001110;
   assign rom_data[11529]=8'b01011111;
   assign rom_data[11530]=8'b01001110;
   assign rom_data[11531]=8'b01100001;
   assign rom_data[11532]=8'b01001110;
   assign rom_data[11533]=8'b01100010;
   assign rom_data[11534]=8'b01001110;
   assign rom_data[11535]=8'b01100011;
   assign rom_data[11536]=8'b01001110;
   assign rom_data[11537]=8'b01100101;
   assign rom_data[11538]=8'b01001101;
   assign rom_data[11539]=8'b01100110;
   assign rom_data[11540]=8'b01001101;
   assign rom_data[11541]=8'b01101000;
   assign rom_data[11542]=8'b01001101;
   assign rom_data[11543]=8'b01101001;
   assign rom_data[11544]=8'b01001101;
   assign rom_data[11545]=8'b01101010;
   assign rom_data[11546]=8'b01001101;
   assign rom_data[11547]=8'b01101100;
   assign rom_data[11548]=8'b01001101;
   assign rom_data[11549]=8'b01101101;
   assign rom_data[11550]=8'b01001101;
   assign rom_data[11551]=8'b01101110;
   assign rom_data[11552]=8'b01001101;
   assign rom_data[11553]=8'b01110000;
   assign rom_data[11554]=8'b01001101;
   assign rom_data[11555]=8'b01110001;
   assign rom_data[11556]=8'b01001101;
   assign rom_data[11557]=8'b01110010;
   assign rom_data[11558]=8'b01001101;
   assign rom_data[11559]=8'b01110100;
   assign rom_data[11560]=8'b01001101;
   assign rom_data[11561]=8'b01110101;
   assign rom_data[11562]=8'b01001101;
   assign rom_data[11563]=8'b01110110;
   assign rom_data[11564]=8'b01001101;
   assign rom_data[11565]=8'b01110111;
   assign rom_data[11566]=8'b01001101;
   assign rom_data[11567]=8'b01111001;
   assign rom_data[11568]=8'b01001101;
   assign rom_data[11569]=8'b01111010;
   assign rom_data[11570]=8'b01001101;
   assign rom_data[11571]=8'b01111011;
   assign rom_data[11572]=8'b01001101;
   assign rom_data[11573]=8'b01111100;
   assign rom_data[11574]=8'b01001101;
   assign rom_data[11575]=8'b01111101;
   assign rom_data[11576]=8'b01001101;
   assign rom_data[11577]=8'b01111110;
   assign rom_data[11578]=8'b01001101;
   assign rom_data[11579]=8'b01111111;
   assign rom_data[11580]=8'b01001101;
   assign rom_data[11581]=8'b10000000;
   assign rom_data[11582]=8'b01001101;
   assign rom_data[11583]=8'b10000001;
   assign rom_data[11584]=8'b01001101;
   assign rom_data[11585]=8'b10000010;
   assign rom_data[11586]=8'b01001101;
   assign rom_data[11587]=8'b10000011;
   assign rom_data[11588]=8'b01001101;
   assign rom_data[11589]=8'b10000100;
   assign rom_data[11590]=8'b01001101;
   assign rom_data[11591]=8'b10000101;
   assign rom_data[11592]=8'b01001101;
   assign rom_data[11593]=8'b10000110;
   assign rom_data[11594]=8'b01001101;
   assign rom_data[11595]=8'b10000110;
   assign rom_data[11596]=8'b01001101;
   assign rom_data[11597]=8'b10000111;
   assign rom_data[11598]=8'b01001101;
   assign rom_data[11599]=8'b10001000;
   assign rom_data[11600]=8'b01001101;
   assign rom_data[11601]=8'b10001000;
   assign rom_data[11602]=8'b01001101;
   assign rom_data[11603]=8'b10001001;
   assign rom_data[11604]=8'b01001101;
   assign rom_data[11605]=8'b10001001;
   assign rom_data[11606]=8'b01001101;
   assign rom_data[11607]=8'b10001001;
   assign rom_data[11608]=8'b01001101;
   assign rom_data[11609]=8'b10001010;
   assign rom_data[11610]=8'b01001100;
   assign rom_data[11611]=8'b10001010;
   assign rom_data[11612]=8'b01001100;
   assign rom_data[11613]=8'b10001010;
   assign rom_data[11614]=8'b01001100;
   assign rom_data[11615]=8'b10001010;
   assign rom_data[11616]=8'b01001100;
   assign rom_data[11617]=8'b10001010;
   assign rom_data[11618]=8'b01001100;
   assign rom_data[11619]=8'b10001001;
   assign rom_data[11620]=8'b01001100;
   assign rom_data[11621]=8'b10001001;
   assign rom_data[11622]=8'b01001100;
   assign rom_data[11623]=8'b10001001;
   assign rom_data[11624]=8'b01001100;
   assign rom_data[11625]=8'b10001000;
   assign rom_data[11626]=8'b01001100;
   assign rom_data[11627]=8'b10001000;
   assign rom_data[11628]=8'b01001100;
   assign rom_data[11629]=8'b10000111;
   assign rom_data[11630]=8'b01001100;
   assign rom_data[11631]=8'b10000111;
   assign rom_data[11632]=8'b01001100;
   assign rom_data[11633]=8'b10000110;
   assign rom_data[11634]=8'b01001100;
   assign rom_data[11635]=8'b10000101;
   assign rom_data[11636]=8'b01001100;
   assign rom_data[11637]=8'b10000100;
   assign rom_data[11638]=8'b01001100;
   assign rom_data[11639]=8'b10000011;
   assign rom_data[11640]=8'b01001100;
   assign rom_data[11641]=8'b10000011;
   assign rom_data[11642]=8'b01001100;
   assign rom_data[11643]=8'b10000010;
   assign rom_data[11644]=8'b01001100;
   assign rom_data[11645]=8'b10000001;
   assign rom_data[11646]=8'b01001100;
   assign rom_data[11647]=8'b10000000;
   assign rom_data[11648]=8'b01001100;
   assign rom_data[11649]=8'b01111110;
   assign rom_data[11650]=8'b01001100;
   assign rom_data[11651]=8'b01111101;
   assign rom_data[11652]=8'b01001100;
   assign rom_data[11653]=8'b01111100;
   assign rom_data[11654]=8'b01001100;
   assign rom_data[11655]=8'b01111011;
   assign rom_data[11656]=8'b01001100;
   assign rom_data[11657]=8'b01111010;
   assign rom_data[11658]=8'b01001100;
   assign rom_data[11659]=8'b01111001;
   assign rom_data[11660]=8'b01001100;
   assign rom_data[11661]=8'b01110111;
   assign rom_data[11662]=8'b01001100;
   assign rom_data[11663]=8'b01110110;
   assign rom_data[11664]=8'b01001100;
   assign rom_data[11665]=8'b01110101;
   assign rom_data[11666]=8'b01001100;
   assign rom_data[11667]=8'b01110100;
   assign rom_data[11668]=8'b01001100;
   assign rom_data[11669]=8'b01110010;
   assign rom_data[11670]=8'b01001100;
   assign rom_data[11671]=8'b01110001;
   assign rom_data[11672]=8'b01001100;
   assign rom_data[11673]=8'b01110000;
   assign rom_data[11674]=8'b01001100;
   assign rom_data[11675]=8'b01101110;
   assign rom_data[11676]=8'b01001100;
   assign rom_data[11677]=8'b01101101;
   assign rom_data[11678]=8'b01001100;
   assign rom_data[11679]=8'b01101100;
   assign rom_data[11680]=8'b01001100;
   assign rom_data[11681]=8'b01101010;
   assign rom_data[11682]=8'b01001011;
   assign rom_data[11683]=8'b01101001;
   assign rom_data[11684]=8'b01001011;
   assign rom_data[11685]=8'b01100111;
   assign rom_data[11686]=8'b01001011;
   assign rom_data[11687]=8'b01100110;
   assign rom_data[11688]=8'b01001011;
   assign rom_data[11689]=8'b01100101;
   assign rom_data[11690]=8'b01001011;
   assign rom_data[11691]=8'b01100011;
   assign rom_data[11692]=8'b01001011;
   assign rom_data[11693]=8'b01100010;
   assign rom_data[11694]=8'b01001011;
   assign rom_data[11695]=8'b01100000;
   assign rom_data[11696]=8'b01001011;
   assign rom_data[11697]=8'b01011111;
   assign rom_data[11698]=8'b01001011;
   assign rom_data[11699]=8'b01011110;
   assign rom_data[11700]=8'b01001011;
   assign rom_data[11701]=8'b01011100;
   assign rom_data[11702]=8'b01001011;
   assign rom_data[11703]=8'b01011011;
   assign rom_data[11704]=8'b01001011;
   assign rom_data[11705]=8'b01011001;
   assign rom_data[11706]=8'b01001011;
   assign rom_data[11707]=8'b01011000;
   assign rom_data[11708]=8'b01001011;
   assign rom_data[11709]=8'b01010111;
   assign rom_data[11710]=8'b01001011;
   assign rom_data[11711]=8'b01010101;
   assign rom_data[11712]=8'b01001011;
   assign rom_data[11713]=8'b01010100;
   assign rom_data[11714]=8'b01001011;
   assign rom_data[11715]=8'b01010010;
   assign rom_data[11716]=8'b01001011;
   assign rom_data[11717]=8'b01010001;
   assign rom_data[11718]=8'b01001011;
   assign rom_data[11719]=8'b01010000;
   assign rom_data[11720]=8'b01001011;
   assign rom_data[11721]=8'b01001110;
   assign rom_data[11722]=8'b01001011;
   assign rom_data[11723]=8'b01001101;
   assign rom_data[11724]=8'b01001011;
   assign rom_data[11725]=8'b01001100;
   assign rom_data[11726]=8'b01001011;
   assign rom_data[11727]=8'b01001010;
   assign rom_data[11728]=8'b01001011;
   assign rom_data[11729]=8'b01001001;
   assign rom_data[11730]=8'b01001011;
   assign rom_data[11731]=8'b01000111;
   assign rom_data[11732]=8'b01001011;
   assign rom_data[11733]=8'b01000110;
   assign rom_data[11734]=8'b01001011;
   assign rom_data[11735]=8'b01000101;
   assign rom_data[11736]=8'b01001011;
   assign rom_data[11737]=8'b01000100;
   assign rom_data[11738]=8'b01001011;
   assign rom_data[11739]=8'b01000010;
   assign rom_data[11740]=8'b01001011;
   assign rom_data[11741]=8'b01000001;
   assign rom_data[11742]=8'b01001011;
   assign rom_data[11743]=8'b01000000;
   assign rom_data[11744]=8'b01001011;
   assign rom_data[11745]=8'b00111110;
   assign rom_data[11746]=8'b01001011;
   assign rom_data[11747]=8'b00111101;
   assign rom_data[11748]=8'b01001011;
   assign rom_data[11749]=8'b00111100;
   assign rom_data[11750]=8'b01001011;
   assign rom_data[11751]=8'b00111011;
   assign rom_data[11752]=8'b01001011;
   assign rom_data[11753]=8'b00111010;
   assign rom_data[11754]=8'b01001011;
   assign rom_data[11755]=8'b00111001;
   assign rom_data[11756]=8'b01001011;
   assign rom_data[11757]=8'b00110111;
   assign rom_data[11758]=8'b01001011;
   assign rom_data[11759]=8'b00110110;
   assign rom_data[11760]=8'b01001011;
   assign rom_data[11761]=8'b00110101;
   assign rom_data[11762]=8'b01001011;
   assign rom_data[11763]=8'b00110100;
   assign rom_data[11764]=8'b01001010;
   assign rom_data[11765]=8'b00110011;
   assign rom_data[11766]=8'b01001010;
   assign rom_data[11767]=8'b00110011;
   assign rom_data[11768]=8'b01001010;
   assign rom_data[11769]=8'b00110010;
   assign rom_data[11770]=8'b01001010;
   assign rom_data[11771]=8'b00110001;
   assign rom_data[11772]=8'b01001010;
   assign rom_data[11773]=8'b00110000;
   assign rom_data[11774]=8'b01001010;
   assign rom_data[11775]=8'b00101111;
   assign rom_data[11776]=8'b01001010;
   assign rom_data[11777]=8'b00101111;
   assign rom_data[11778]=8'b01001010;
   assign rom_data[11779]=8'b00101110;
   assign rom_data[11780]=8'b01001010;
   assign rom_data[11781]=8'b00101110;
   assign rom_data[11782]=8'b01001010;
   assign rom_data[11783]=8'b00101101;
   assign rom_data[11784]=8'b01001010;
   assign rom_data[11785]=8'b00101101;
   assign rom_data[11786]=8'b01001010;
   assign rom_data[11787]=8'b00101100;
   assign rom_data[11788]=8'b01001010;
   assign rom_data[11789]=8'b00101100;
   assign rom_data[11790]=8'b01001010;
   assign rom_data[11791]=8'b00101100;
   assign rom_data[11792]=8'b01001010;
   assign rom_data[11793]=8'b00101100;
   assign rom_data[11794]=8'b01001010;
   assign rom_data[11795]=8'b00101100;
   assign rom_data[11796]=8'b01001010;
   assign rom_data[11797]=8'b00101100;
   assign rom_data[11798]=8'b01001010;
   assign rom_data[11799]=8'b00101100;
   assign rom_data[11800]=8'b01001010;
   assign rom_data[11801]=8'b00101101;
   assign rom_data[11802]=8'b01001010;
   assign rom_data[11803]=8'b00101101;
   assign rom_data[11804]=8'b01001010;
   assign rom_data[11805]=8'b00101101;
   assign rom_data[11806]=8'b01001010;
   assign rom_data[11807]=8'b00101110;
   assign rom_data[11808]=8'b01001010;
   assign rom_data[11809]=8'b00101111;
   assign rom_data[11810]=8'b01001010;
   assign rom_data[11811]=8'b00101111;
   assign rom_data[11812]=8'b01001010;
   assign rom_data[11813]=8'b00110000;
   assign rom_data[11814]=8'b01001010;
   assign rom_data[11815]=8'b00110001;
   assign rom_data[11816]=8'b01001010;
   assign rom_data[11817]=8'b00110010;
   assign rom_data[11818]=8'b01001010;
   assign rom_data[11819]=8'b00110010;
   assign rom_data[11820]=8'b01001010;
   assign rom_data[11821]=8'b00110011;
   assign rom_data[11822]=8'b01001010;
   assign rom_data[11823]=8'b00110100;
   assign rom_data[11824]=8'b01001010;
   assign rom_data[11825]=8'b00110101;
   assign rom_data[11826]=8'b01001010;
   assign rom_data[11827]=8'b00110110;
   assign rom_data[11828]=8'b01001010;
   assign rom_data[11829]=8'b00110111;
   assign rom_data[11830]=8'b01001001;
   assign rom_data[11831]=8'b00111001;
   assign rom_data[11832]=8'b01001001;
   assign rom_data[11833]=8'b00111010;
   assign rom_data[11834]=8'b01001001;
   assign rom_data[11835]=8'b00111011;
   assign rom_data[11836]=8'b01001001;
   assign rom_data[11837]=8'b00111100;
   assign rom_data[11838]=8'b01001001;
   assign rom_data[11839]=8'b00111101;
   assign rom_data[11840]=8'b01001001;
   assign rom_data[11841]=8'b00111110;
   assign rom_data[11842]=8'b01001001;
   assign rom_data[11843]=8'b01000000;
   assign rom_data[11844]=8'b01001001;
   assign rom_data[11845]=8'b01000001;
   assign rom_data[11846]=8'b01001001;
   assign rom_data[11847]=8'b01000010;
   assign rom_data[11848]=8'b01001001;
   assign rom_data[11849]=8'b01000100;
   assign rom_data[11850]=8'b01001001;
   assign rom_data[11851]=8'b01000101;
   assign rom_data[11852]=8'b01001001;
   assign rom_data[11853]=8'b01000110;
   assign rom_data[11854]=8'b01001001;
   assign rom_data[11855]=8'b01001000;
   assign rom_data[11856]=8'b01001001;
   assign rom_data[11857]=8'b01001001;
   assign rom_data[11858]=8'b01001001;
   assign rom_data[11859]=8'b01001010;
   assign rom_data[11860]=8'b01001001;
   assign rom_data[11861]=8'b01001100;
   assign rom_data[11862]=8'b01001001;
   assign rom_data[11863]=8'b01001101;
   assign rom_data[11864]=8'b01001001;
   assign rom_data[11865]=8'b01001110;
   assign rom_data[11866]=8'b01001001;
   assign rom_data[11867]=8'b01010000;
   assign rom_data[11868]=8'b01001001;
   assign rom_data[11869]=8'b01010001;
   assign rom_data[11870]=8'b01001001;
   assign rom_data[11871]=8'b01010011;
   assign rom_data[11872]=8'b01001001;
   assign rom_data[11873]=8'b01010100;
   assign rom_data[11874]=8'b01001001;
   assign rom_data[11875]=8'b01010101;
   assign rom_data[11876]=8'b01001001;
   assign rom_data[11877]=8'b01010111;
   assign rom_data[11878]=8'b01001001;
   assign rom_data[11879]=8'b01011000;
   assign rom_data[11880]=8'b01001001;
   assign rom_data[11881]=8'b01011010;
   assign rom_data[11882]=8'b01001001;
   assign rom_data[11883]=8'b01011011;
   assign rom_data[11884]=8'b01001001;
   assign rom_data[11885]=8'b01011100;
   assign rom_data[11886]=8'b01001001;
   assign rom_data[11887]=8'b01011110;
   assign rom_data[11888]=8'b01001001;
   assign rom_data[11889]=8'b01011111;
   assign rom_data[11890]=8'b01001001;
   assign rom_data[11891]=8'b01100001;
   assign rom_data[11892]=8'b01001001;
   assign rom_data[11893]=8'b01100010;
   assign rom_data[11894]=8'b01001001;
   assign rom_data[11895]=8'b01100011;
   assign rom_data[11896]=8'b01001001;
   assign rom_data[11897]=8'b01100101;
   assign rom_data[11898]=8'b01001001;
   assign rom_data[11899]=8'b01100110;
   assign rom_data[11900]=8'b01001001;
   assign rom_data[11901]=8'b01101000;
   assign rom_data[11902]=8'b01001001;
   assign rom_data[11903]=8'b01101001;
   assign rom_data[11904]=8'b01001001;
   assign rom_data[11905]=8'b01101010;
   assign rom_data[11906]=8'b01001001;
   assign rom_data[11907]=8'b01101100;
   assign rom_data[11908]=8'b01001001;
   assign rom_data[11909]=8'b01101101;
   assign rom_data[11910]=8'b01001001;
   assign rom_data[11911]=8'b01101110;
   assign rom_data[11912]=8'b01001001;
   assign rom_data[11913]=8'b01110000;
   assign rom_data[11914]=8'b01001000;
   assign rom_data[11915]=8'b01110001;
   assign rom_data[11916]=8'b01001000;
   assign rom_data[11917]=8'b01110010;
   assign rom_data[11918]=8'b01001000;
   assign rom_data[11919]=8'b01110100;
   assign rom_data[11920]=8'b01001000;
   assign rom_data[11921]=8'b01110101;
   assign rom_data[11922]=8'b01001000;
   assign rom_data[11923]=8'b01110110;
   assign rom_data[11924]=8'b01001000;
   assign rom_data[11925]=8'b01110111;
   assign rom_data[11926]=8'b01001000;
   assign rom_data[11927]=8'b01111001;
   assign rom_data[11928]=8'b01001000;
   assign rom_data[11929]=8'b01111010;
   assign rom_data[11930]=8'b01001000;
   assign rom_data[11931]=8'b01111011;
   assign rom_data[11932]=8'b01001000;
   assign rom_data[11933]=8'b01111100;
   assign rom_data[11934]=8'b01001000;
   assign rom_data[11935]=8'b01111101;
   assign rom_data[11936]=8'b01001000;
   assign rom_data[11937]=8'b01111110;
   assign rom_data[11938]=8'b01001000;
   assign rom_data[11939]=8'b01111111;
   assign rom_data[11940]=8'b01001000;
   assign rom_data[11941]=8'b10000000;
   assign rom_data[11942]=8'b01001000;
   assign rom_data[11943]=8'b10000001;
   assign rom_data[11944]=8'b01001000;
   assign rom_data[11945]=8'b10000010;
   assign rom_data[11946]=8'b01001000;
   assign rom_data[11947]=8'b10000011;
   assign rom_data[11948]=8'b01001000;
   assign rom_data[11949]=8'b10000100;
   assign rom_data[11950]=8'b01001000;
   assign rom_data[11951]=8'b10000101;
   assign rom_data[11952]=8'b01001000;
   assign rom_data[11953]=8'b10000110;
   assign rom_data[11954]=8'b01001000;
   assign rom_data[11955]=8'b10000110;
   assign rom_data[11956]=8'b01001000;
   assign rom_data[11957]=8'b10000111;
   assign rom_data[11958]=8'b01001000;
   assign rom_data[11959]=8'b10001000;
   assign rom_data[11960]=8'b01001000;
   assign rom_data[11961]=8'b10001000;
   assign rom_data[11962]=8'b01001000;
   assign rom_data[11963]=8'b10001001;
   assign rom_data[11964]=8'b01001000;
   assign rom_data[11965]=8'b10001001;
   assign rom_data[11966]=8'b01001000;
   assign rom_data[11967]=8'b10001001;
   assign rom_data[11968]=8'b01001000;
   assign rom_data[11969]=8'b10001010;
   assign rom_data[11970]=8'b01001000;
   assign rom_data[11971]=8'b10001010;
   assign rom_data[11972]=8'b01001000;
   assign rom_data[11973]=8'b10001010;
   assign rom_data[11974]=8'b01001000;
   assign rom_data[11975]=8'b10001010;
   assign rom_data[11976]=8'b01001000;
   assign rom_data[11977]=8'b10001010;
   assign rom_data[11978]=8'b01001000;
   assign rom_data[11979]=8'b10001001;
   assign rom_data[11980]=8'b01001000;
   assign rom_data[11981]=8'b10001001;
   assign rom_data[11982]=8'b01000111;
   assign rom_data[11983]=8'b10001001;
   assign rom_data[11984]=8'b01000111;
   assign rom_data[11985]=8'b10001000;
   assign rom_data[11986]=8'b01000111;
   assign rom_data[11987]=8'b10001000;
   assign rom_data[11988]=8'b01000111;
   assign rom_data[11989]=8'b10000111;
   assign rom_data[11990]=8'b01000111;
   assign rom_data[11991]=8'b10000111;
   assign rom_data[11992]=8'b01000111;
   assign rom_data[11993]=8'b10000110;
   assign rom_data[11994]=8'b01000111;
   assign rom_data[11995]=8'b10000101;
   assign rom_data[11996]=8'b01000111;
   assign rom_data[11997]=8'b10000100;
   assign rom_data[11998]=8'b01000111;
   assign rom_data[11999]=8'b10000011;
   assign rom_data[12000]=8'b01000111;
   assign rom_data[12001]=8'b10000011;
   assign rom_data[12002]=8'b01000111;
   assign rom_data[12003]=8'b10000010;
   assign rom_data[12004]=8'b01000111;
   assign rom_data[12005]=8'b10000001;
   assign rom_data[12006]=8'b01000111;
   assign rom_data[12007]=8'b01111111;
   assign rom_data[12008]=8'b01000111;
   assign rom_data[12009]=8'b01111110;
   assign rom_data[12010]=8'b01000111;
   assign rom_data[12011]=8'b01111101;
   assign rom_data[12012]=8'b01000111;
   assign rom_data[12013]=8'b01111100;
   assign rom_data[12014]=8'b01000111;
   assign rom_data[12015]=8'b01111011;
   assign rom_data[12016]=8'b01000111;
   assign rom_data[12017]=8'b01111010;
   assign rom_data[12018]=8'b01000111;
   assign rom_data[12019]=8'b01111001;
   assign rom_data[12020]=8'b01000111;
   assign rom_data[12021]=8'b01110111;
   assign rom_data[12022]=8'b01000111;
   assign rom_data[12023]=8'b01110110;
   assign rom_data[12024]=8'b01000111;
   assign rom_data[12025]=8'b01110101;
   assign rom_data[12026]=8'b01000111;
   assign rom_data[12027]=8'b01110100;
   assign rom_data[12028]=8'b01000111;
   assign rom_data[12029]=8'b01110010;
   assign rom_data[12030]=8'b01000111;
   assign rom_data[12031]=8'b01110001;
   assign rom_data[12032]=8'b01000111;
   assign rom_data[12033]=8'b01110000;
   assign rom_data[12034]=8'b01000111;
   assign rom_data[12035]=8'b01101110;
   assign rom_data[12036]=8'b01000111;
   assign rom_data[12037]=8'b01101101;
   assign rom_data[12038]=8'b01000111;
   assign rom_data[12039]=8'b01101100;
   assign rom_data[12040]=8'b01000111;
   assign rom_data[12041]=8'b01101010;
   assign rom_data[12042]=8'b01000111;
   assign rom_data[12043]=8'b01101001;
   assign rom_data[12044]=8'b01000111;
   assign rom_data[12045]=8'b01100111;
   assign rom_data[12046]=8'b01000111;
   assign rom_data[12047]=8'b01100110;
   assign rom_data[12048]=8'b01000111;
   assign rom_data[12049]=8'b01100101;
   assign rom_data[12050]=8'b01000111;
   assign rom_data[12051]=8'b01100011;
   assign rom_data[12052]=8'b01000111;
   assign rom_data[12053]=8'b01100010;
   assign rom_data[12054]=8'b01000111;
   assign rom_data[12055]=8'b01100000;
   assign rom_data[12056]=8'b01000111;
   assign rom_data[12057]=8'b01011111;
   assign rom_data[12058]=8'b01000111;
   assign rom_data[12059]=8'b01011110;
   assign rom_data[12060]=8'b01000110;
   assign rom_data[12061]=8'b01011100;
   assign rom_data[12062]=8'b01000110;
   assign rom_data[12063]=8'b01011011;
   assign rom_data[12064]=8'b01000110;
   assign rom_data[12065]=8'b01011001;
   assign rom_data[12066]=8'b01000110;
   assign rom_data[12067]=8'b01011000;
   assign rom_data[12068]=8'b01000110;
   assign rom_data[12069]=8'b01010111;
   assign rom_data[12070]=8'b01000110;
   assign rom_data[12071]=8'b01010101;
   assign rom_data[12072]=8'b01000110;
   assign rom_data[12073]=8'b01010100;
   assign rom_data[12074]=8'b01000110;
   assign rom_data[12075]=8'b01010010;
   assign rom_data[12076]=8'b01000110;
   assign rom_data[12077]=8'b01010001;
   assign rom_data[12078]=8'b01000110;
   assign rom_data[12079]=8'b01010000;
   assign rom_data[12080]=8'b01000110;
   assign rom_data[12081]=8'b01001110;
   assign rom_data[12082]=8'b01000110;
   assign rom_data[12083]=8'b01001101;
   assign rom_data[12084]=8'b01000110;
   assign rom_data[12085]=8'b01001100;
   assign rom_data[12086]=8'b01000110;
   assign rom_data[12087]=8'b01001010;
   assign rom_data[12088]=8'b01000110;
   assign rom_data[12089]=8'b01001001;
   assign rom_data[12090]=8'b01000110;
   assign rom_data[12091]=8'b01000111;
   assign rom_data[12092]=8'b01000110;
   assign rom_data[12093]=8'b01000110;
   assign rom_data[12094]=8'b01000110;
   assign rom_data[12095]=8'b01000101;
   assign rom_data[12096]=8'b01000110;
   assign rom_data[12097]=8'b01000100;
   assign rom_data[12098]=8'b01000110;
   assign rom_data[12099]=8'b01000010;
   assign rom_data[12100]=8'b01000110;
   assign rom_data[12101]=8'b01000001;
   assign rom_data[12102]=8'b01000110;
   assign rom_data[12103]=8'b01000000;
   assign rom_data[12104]=8'b01000110;
   assign rom_data[12105]=8'b00111110;
   assign rom_data[12106]=8'b01000110;
   assign rom_data[12107]=8'b00111101;
   assign rom_data[12108]=8'b01000110;
   assign rom_data[12109]=8'b00111100;
   assign rom_data[12110]=8'b01000110;
   assign rom_data[12111]=8'b00111011;
   assign rom_data[12112]=8'b01000110;
   assign rom_data[12113]=8'b00111010;
   assign rom_data[12114]=8'b01000110;
   assign rom_data[12115]=8'b00111001;
   assign rom_data[12116]=8'b01000110;
   assign rom_data[12117]=8'b00110111;
   assign rom_data[12118]=8'b01000110;
   assign rom_data[12119]=8'b00110110;
   assign rom_data[12120]=8'b01000110;
   assign rom_data[12121]=8'b00110101;
   assign rom_data[12122]=8'b01000110;
   assign rom_data[12123]=8'b00110100;
   assign rom_data[12124]=8'b01000110;
   assign rom_data[12125]=8'b00110011;
   assign rom_data[12126]=8'b01000110;
   assign rom_data[12127]=8'b00110011;
   assign rom_data[12128]=8'b01000110;
   assign rom_data[12129]=8'b00110010;
   assign rom_data[12130]=8'b01000110;
   assign rom_data[12131]=8'b00110001;
   assign rom_data[12132]=8'b01000110;
   assign rom_data[12133]=8'b00110000;
   assign rom_data[12134]=8'b01000110;
   assign rom_data[12135]=8'b00101111;
   assign rom_data[12136]=8'b01000101;
   assign rom_data[12137]=8'b00101111;
   assign rom_data[12138]=8'b01000101;
   assign rom_data[12139]=8'b00101110;
   assign rom_data[12140]=8'b01000101;
   assign rom_data[12141]=8'b00101110;
   assign rom_data[12142]=8'b01000101;
   assign rom_data[12143]=8'b00101101;
   assign rom_data[12144]=8'b01000101;
   assign rom_data[12145]=8'b00101101;
   assign rom_data[12146]=8'b01000101;
   assign rom_data[12147]=8'b00101100;
   assign rom_data[12148]=8'b01000101;
   assign rom_data[12149]=8'b00101100;
   assign rom_data[12150]=8'b01000101;
   assign rom_data[12151]=8'b00101100;
   assign rom_data[12152]=8'b01000101;
   assign rom_data[12153]=8'b00101100;
   assign rom_data[12154]=8'b01000101;
   assign rom_data[12155]=8'b00101100;
   assign rom_data[12156]=8'b01000101;
   assign rom_data[12157]=8'b00101100;
   assign rom_data[12158]=8'b01000101;
   assign rom_data[12159]=8'b00101100;
   assign rom_data[12160]=8'b01000101;
   assign rom_data[12161]=8'b00101101;
   assign rom_data[12162]=8'b01000101;
   assign rom_data[12163]=8'b00101101;
   assign rom_data[12164]=8'b01000101;
   assign rom_data[12165]=8'b00101101;
   assign rom_data[12166]=8'b01000101;
   assign rom_data[12167]=8'b00101110;
   assign rom_data[12168]=8'b01000101;
   assign rom_data[12169]=8'b00101111;
   assign rom_data[12170]=8'b01000101;
   assign rom_data[12171]=8'b00101111;
   assign rom_data[12172]=8'b01000101;
   assign rom_data[12173]=8'b00110000;
   assign rom_data[12174]=8'b01000101;
   assign rom_data[12175]=8'b00110001;
   assign rom_data[12176]=8'b01000101;
   assign rom_data[12177]=8'b00110010;
   assign rom_data[12178]=8'b01000101;
   assign rom_data[12179]=8'b00110010;
   assign rom_data[12180]=8'b01000101;
   assign rom_data[12181]=8'b00110011;
   assign rom_data[12182]=8'b01000101;
   assign rom_data[12183]=8'b00110100;
   assign rom_data[12184]=8'b01000101;
   assign rom_data[12185]=8'b00110101;
   assign rom_data[12186]=8'b01000101;
   assign rom_data[12187]=8'b00110110;
   assign rom_data[12188]=8'b01000101;
   assign rom_data[12189]=8'b00110111;
   assign rom_data[12190]=8'b01000101;
   assign rom_data[12191]=8'b00111001;
   assign rom_data[12192]=8'b01000101;
   assign rom_data[12193]=8'b00111010;
   assign rom_data[12194]=8'b01000101;
   assign rom_data[12195]=8'b00111011;
   assign rom_data[12196]=8'b01000101;
   assign rom_data[12197]=8'b00111100;
   assign rom_data[12198]=8'b01000101;
   assign rom_data[12199]=8'b00111101;
   assign rom_data[12200]=8'b01000101;
   assign rom_data[12201]=8'b00111110;
   assign rom_data[12202]=8'b01000101;
   assign rom_data[12203]=8'b01000000;
   assign rom_data[12204]=8'b01000101;
   assign rom_data[12205]=8'b01000001;
   assign rom_data[12206]=8'b01000100;
   assign rom_data[12207]=8'b01000010;
   assign rom_data[12208]=8'b01000100;
   assign rom_data[12209]=8'b01000100;
   assign rom_data[12210]=8'b01000100;
   assign rom_data[12211]=8'b01000101;
   assign rom_data[12212]=8'b01000100;
   assign rom_data[12213]=8'b01000110;
   assign rom_data[12214]=8'b01000100;
   assign rom_data[12215]=8'b01001000;
   assign rom_data[12216]=8'b01000100;
   assign rom_data[12217]=8'b01001001;
   assign rom_data[12218]=8'b01000100;
   assign rom_data[12219]=8'b01001010;
   assign rom_data[12220]=8'b01000100;
   assign rom_data[12221]=8'b01001100;
   assign rom_data[12222]=8'b01000100;
   assign rom_data[12223]=8'b01001101;
   assign rom_data[12224]=8'b01000100;
   assign rom_data[12225]=8'b01001110;
   assign rom_data[12226]=8'b01000100;
   assign rom_data[12227]=8'b01010000;
   assign rom_data[12228]=8'b01000100;
   assign rom_data[12229]=8'b01010001;
   assign rom_data[12230]=8'b01000100;
   assign rom_data[12231]=8'b01010011;
   assign rom_data[12232]=8'b01000100;
   assign rom_data[12233]=8'b01010100;
   assign rom_data[12234]=8'b01000100;
   assign rom_data[12235]=8'b01010101;
   assign rom_data[12236]=8'b01000100;
   assign rom_data[12237]=8'b01010111;
   assign rom_data[12238]=8'b01000100;
   assign rom_data[12239]=8'b01011000;
   assign rom_data[12240]=8'b01000100;
   assign rom_data[12241]=8'b01011010;
   assign rom_data[12242]=8'b01000100;
   assign rom_data[12243]=8'b01011011;
   assign rom_data[12244]=8'b01000100;
   assign rom_data[12245]=8'b01011100;
   assign rom_data[12246]=8'b01000100;
   assign rom_data[12247]=8'b01011110;
   assign rom_data[12248]=8'b01000100;
   assign rom_data[12249]=8'b01011111;
   assign rom_data[12250]=8'b01000100;
   assign rom_data[12251]=8'b01100001;
   assign rom_data[12252]=8'b01000100;
   assign rom_data[12253]=8'b01100010;
   assign rom_data[12254]=8'b01000100;
   assign rom_data[12255]=8'b01100011;
   assign rom_data[12256]=8'b01000100;
   assign rom_data[12257]=8'b01100101;
   assign rom_data[12258]=8'b01000100;
   assign rom_data[12259]=8'b01100110;
   assign rom_data[12260]=8'b01000100;
   assign rom_data[12261]=8'b01101000;
   assign rom_data[12262]=8'b01000100;
   assign rom_data[12263]=8'b01101001;
   assign rom_data[12264]=8'b01000100;
   assign rom_data[12265]=8'b01101010;
   assign rom_data[12266]=8'b01000100;
   assign rom_data[12267]=8'b01101100;
   assign rom_data[12268]=8'b01000100;
   assign rom_data[12269]=8'b01101101;
   assign rom_data[12270]=8'b01000100;
   assign rom_data[12271]=8'b01101110;
   assign rom_data[12272]=8'b01000100;
   assign rom_data[12273]=8'b01110000;
   assign rom_data[12274]=8'b01000100;
   assign rom_data[12275]=8'b01110001;
   assign rom_data[12276]=8'b01000100;
   assign rom_data[12277]=8'b01110010;
   assign rom_data[12278]=8'b01000100;
   assign rom_data[12279]=8'b01110100;
   assign rom_data[12280]=8'b01000100;
   assign rom_data[12281]=8'b01110101;
   assign rom_data[12282]=8'b01000100;
   assign rom_data[12283]=8'b01110110;
   assign rom_data[12284]=8'b01000100;
   assign rom_data[12285]=8'b01110111;
   assign rom_data[12286]=8'b01000100;
   assign rom_data[12287]=8'b01111001;
   assign rom_data[12288]=8'b01000011;
   assign rom_data[12289]=8'b01111010;
   assign rom_data[12290]=8'b01000011;
   assign rom_data[12291]=8'b01111011;
   assign rom_data[12292]=8'b01000011;
   assign rom_data[12293]=8'b01111100;
   assign rom_data[12294]=8'b01000011;
   assign rom_data[12295]=8'b01111101;
   assign rom_data[12296]=8'b01000011;
   assign rom_data[12297]=8'b01111110;
   assign rom_data[12298]=8'b01000011;
   assign rom_data[12299]=8'b01111111;
   assign rom_data[12300]=8'b01000011;
   assign rom_data[12301]=8'b10000000;
   assign rom_data[12302]=8'b01000011;
   assign rom_data[12303]=8'b10000001;
   assign rom_data[12304]=8'b01000011;
   assign rom_data[12305]=8'b10000010;
   assign rom_data[12306]=8'b01000011;
   assign rom_data[12307]=8'b10000011;
   assign rom_data[12308]=8'b01000011;
   assign rom_data[12309]=8'b10000100;
   assign rom_data[12310]=8'b01000011;
   assign rom_data[12311]=8'b10000101;
   assign rom_data[12312]=8'b01000011;
   assign rom_data[12313]=8'b10000110;
   assign rom_data[12314]=8'b01000011;
   assign rom_data[12315]=8'b10000110;
   assign rom_data[12316]=8'b01000011;
   assign rom_data[12317]=8'b10000111;
   assign rom_data[12318]=8'b01000011;
   assign rom_data[12319]=8'b10001000;
   assign rom_data[12320]=8'b01000011;
   assign rom_data[12321]=8'b10001000;
   assign rom_data[12322]=8'b01000011;
   assign rom_data[12323]=8'b10001001;
   assign rom_data[12324]=8'b01000011;
   assign rom_data[12325]=8'b10001001;
   assign rom_data[12326]=8'b01000011;
   assign rom_data[12327]=8'b10001001;
   assign rom_data[12328]=8'b01000011;
   assign rom_data[12329]=8'b10001010;
   assign rom_data[12330]=8'b01000011;
   assign rom_data[12331]=8'b10001010;
   assign rom_data[12332]=8'b01000011;
   assign rom_data[12333]=8'b10001010;
   assign rom_data[12334]=8'b01000011;
   assign rom_data[12335]=8'b10001010;
   assign rom_data[12336]=8'b01000011;
   assign rom_data[12337]=8'b10001010;
   assign rom_data[12338]=8'b01000011;
   assign rom_data[12339]=8'b10001001;
   assign rom_data[12340]=8'b01000011;
   assign rom_data[12341]=8'b10001001;
   assign rom_data[12342]=8'b01000011;
   assign rom_data[12343]=8'b10001001;
   assign rom_data[12344]=8'b01000011;
   assign rom_data[12345]=8'b10001000;
   assign rom_data[12346]=8'b01000011;
   assign rom_data[12347]=8'b10001000;
   assign rom_data[12348]=8'b01000011;
   assign rom_data[12349]=8'b10000111;
   assign rom_data[12350]=8'b01000011;
   assign rom_data[12351]=8'b10000111;
   assign rom_data[12352]=8'b01000011;
   assign rom_data[12353]=8'b10000110;
   assign rom_data[12354]=8'b01000010;
   assign rom_data[12355]=8'b10000101;
   assign rom_data[12356]=8'b01000010;
   assign rom_data[12357]=8'b10000100;
   assign rom_data[12358]=8'b01000010;
   assign rom_data[12359]=8'b10000011;
   assign rom_data[12360]=8'b01000010;
   assign rom_data[12361]=8'b10000011;
   assign rom_data[12362]=8'b01000010;
   assign rom_data[12363]=8'b10000010;
   assign rom_data[12364]=8'b01000010;
   assign rom_data[12365]=8'b10000001;
   assign rom_data[12366]=8'b01000010;
   assign rom_data[12367]=8'b01111111;
   assign rom_data[12368]=8'b01000010;
   assign rom_data[12369]=8'b01111110;
   assign rom_data[12370]=8'b01000010;
   assign rom_data[12371]=8'b01111101;
   assign rom_data[12372]=8'b01000010;
   assign rom_data[12373]=8'b01111100;
   assign rom_data[12374]=8'b01000010;
   assign rom_data[12375]=8'b01111011;
   assign rom_data[12376]=8'b01000010;
   assign rom_data[12377]=8'b01111010;
   assign rom_data[12378]=8'b01000010;
   assign rom_data[12379]=8'b01111001;
   assign rom_data[12380]=8'b01000010;
   assign rom_data[12381]=8'b01110111;
   assign rom_data[12382]=8'b01000010;
   assign rom_data[12383]=8'b01110110;
   assign rom_data[12384]=8'b01000010;
   assign rom_data[12385]=8'b01110101;
   assign rom_data[12386]=8'b01000010;
   assign rom_data[12387]=8'b01110100;
   assign rom_data[12388]=8'b01000010;
   assign rom_data[12389]=8'b01110010;
   assign rom_data[12390]=8'b01000010;
   assign rom_data[12391]=8'b01110001;
   assign rom_data[12392]=8'b01000010;
   assign rom_data[12393]=8'b01110000;
   assign rom_data[12394]=8'b01000010;
   assign rom_data[12395]=8'b01101110;
   assign rom_data[12396]=8'b01000010;
   assign rom_data[12397]=8'b01101101;
   assign rom_data[12398]=8'b01000010;
   assign rom_data[12399]=8'b01101100;
   assign rom_data[12400]=8'b01000010;
   assign rom_data[12401]=8'b01101010;
   assign rom_data[12402]=8'b01000010;
   assign rom_data[12403]=8'b01101001;
   assign rom_data[12404]=8'b01000010;
   assign rom_data[12405]=8'b01100111;
   assign rom_data[12406]=8'b01000010;
   assign rom_data[12407]=8'b01100110;
   assign rom_data[12408]=8'b01000010;
   assign rom_data[12409]=8'b01100101;
   assign rom_data[12410]=8'b01000010;
   assign rom_data[12411]=8'b01100011;
   assign rom_data[12412]=8'b01000010;
   assign rom_data[12413]=8'b01100010;
   assign rom_data[12414]=8'b01000010;
   assign rom_data[12415]=8'b01100000;
   assign rom_data[12416]=8'b01000010;
   assign rom_data[12417]=8'b01011111;
   assign rom_data[12418]=8'b01000010;
   assign rom_data[12419]=8'b01011110;
   assign rom_data[12420]=8'b01000010;
   assign rom_data[12421]=8'b01011100;
   assign rom_data[12422]=8'b01000010;
   assign rom_data[12423]=8'b01011011;
   assign rom_data[12424]=8'b01000010;
   assign rom_data[12425]=8'b01011001;
   assign rom_data[12426]=8'b01000010;
   assign rom_data[12427]=8'b01011000;
   assign rom_data[12428]=8'b01000010;
   assign rom_data[12429]=8'b01010111;
   assign rom_data[12430]=8'b01000010;
   assign rom_data[12431]=8'b01010101;
   assign rom_data[12432]=8'b01000010;
   assign rom_data[12433]=8'b01010100;
   assign rom_data[12434]=8'b01000010;
   assign rom_data[12435]=8'b01010010;
   assign rom_data[12436]=8'b01000001;
   assign rom_data[12437]=8'b01010001;
   assign rom_data[12438]=8'b01000001;
   assign rom_data[12439]=8'b01010000;
   assign rom_data[12440]=8'b01000001;
   assign rom_data[12441]=8'b01001110;
   assign rom_data[12442]=8'b01000001;
   assign rom_data[12443]=8'b01001101;
   assign rom_data[12444]=8'b01000001;
   assign rom_data[12445]=8'b01001100;
   assign rom_data[12446]=8'b01000001;
   assign rom_data[12447]=8'b01001010;
   assign rom_data[12448]=8'b01000001;
   assign rom_data[12449]=8'b01001001;
   assign rom_data[12450]=8'b01000001;
   assign rom_data[12451]=8'b01000111;
   assign rom_data[12452]=8'b01000001;
   assign rom_data[12453]=8'b01000110;
   assign rom_data[12454]=8'b01000001;
   assign rom_data[12455]=8'b01000101;
   assign rom_data[12456]=8'b01000001;
   assign rom_data[12457]=8'b01000100;
   assign rom_data[12458]=8'b01000001;
   assign rom_data[12459]=8'b01000010;
   assign rom_data[12460]=8'b01000001;
   assign rom_data[12461]=8'b01000001;
   assign rom_data[12462]=8'b01000001;
   assign rom_data[12463]=8'b01000000;
   assign rom_data[12464]=8'b01000001;
   assign rom_data[12465]=8'b00111110;
   assign rom_data[12466]=8'b01000001;
   assign rom_data[12467]=8'b00111101;
   assign rom_data[12468]=8'b01000001;
   assign rom_data[12469]=8'b00111100;
   assign rom_data[12470]=8'b01000001;
   assign rom_data[12471]=8'b00111011;
   assign rom_data[12472]=8'b01000001;
   assign rom_data[12473]=8'b00111010;
   assign rom_data[12474]=8'b01000001;
   assign rom_data[12475]=8'b00111001;
   assign rom_data[12476]=8'b01000001;
   assign rom_data[12477]=8'b00110111;
   assign rom_data[12478]=8'b01000001;
   assign rom_data[12479]=8'b00110110;
   assign rom_data[12480]=8'b01000001;
   assign rom_data[12481]=8'b00110101;
   assign rom_data[12482]=8'b01000001;
   assign rom_data[12483]=8'b00110100;
   assign rom_data[12484]=8'b01000001;
   assign rom_data[12485]=8'b00110011;
   assign rom_data[12486]=8'b01000001;
   assign rom_data[12487]=8'b00110011;
   assign rom_data[12488]=8'b01000001;
   assign rom_data[12489]=8'b00110010;
   assign rom_data[12490]=8'b01000001;
   assign rom_data[12491]=8'b00110001;
   assign rom_data[12492]=8'b01000001;
   assign rom_data[12493]=8'b00110000;
   assign rom_data[12494]=8'b01000001;
   assign rom_data[12495]=8'b00101111;
   assign rom_data[12496]=8'b01000001;
   assign rom_data[12497]=8'b00101111;
   assign rom_data[12498]=8'b01000001;
   assign rom_data[12499]=8'b00101110;
   assign rom_data[12500]=8'b01000001;
   assign rom_data[12501]=8'b00101110;
   assign rom_data[12502]=8'b01000001;
   assign rom_data[12503]=8'b00101101;
   assign rom_data[12504]=8'b01000001;
   assign rom_data[12505]=8'b00101101;
   assign rom_data[12506]=8'b01000001;
   assign rom_data[12507]=8'b00101100;
   assign rom_data[12508]=8'b01000000;
   assign rom_data[12509]=8'b00101100;
   assign rom_data[12510]=8'b01000000;
   assign rom_data[12511]=8'b00101100;
   assign rom_data[12512]=8'b01000000;
   assign rom_data[12513]=8'b00101100;
   assign rom_data[12514]=8'b01000000;
   assign rom_data[12515]=8'b00101100;
   assign rom_data[12516]=8'b01000000;
   assign rom_data[12517]=8'b00101100;
   assign rom_data[12518]=8'b01000000;
   assign rom_data[12519]=8'b00101100;
   assign rom_data[12520]=8'b01000000;
   assign rom_data[12521]=8'b00101101;
   assign rom_data[12522]=8'b01000000;
   assign rom_data[12523]=8'b00101101;
   assign rom_data[12524]=8'b01000000;
   assign rom_data[12525]=8'b00101101;
   assign rom_data[12526]=8'b01000000;
   assign rom_data[12527]=8'b00101110;
   assign rom_data[12528]=8'b01000000;
   assign rom_data[12529]=8'b00101111;
   assign rom_data[12530]=8'b01000000;
   assign rom_data[12531]=8'b00101111;
   assign rom_data[12532]=8'b01000000;
   assign rom_data[12533]=8'b00110000;
   assign rom_data[12534]=8'b01000000;
   assign rom_data[12535]=8'b00110001;
   assign rom_data[12536]=8'b01000000;
   assign rom_data[12537]=8'b00110010;
   assign rom_data[12538]=8'b01000000;
   assign rom_data[12539]=8'b00110010;
   assign rom_data[12540]=8'b01000000;
   assign rom_data[12541]=8'b00110011;
   assign rom_data[12542]=8'b01000000;
   assign rom_data[12543]=8'b00110100;
   assign rom_data[12544]=8'b01000000;
   assign rom_data[12545]=8'b00110101;
   assign rom_data[12546]=8'b01000000;
   assign rom_data[12547]=8'b00110110;
   assign rom_data[12548]=8'b01000000;
   assign rom_data[12549]=8'b00110111;
   assign rom_data[12550]=8'b01000000;
   assign rom_data[12551]=8'b00111001;
   assign rom_data[12552]=8'b01000000;
   assign rom_data[12553]=8'b00111010;
   assign rom_data[12554]=8'b01000000;
   assign rom_data[12555]=8'b00111011;
   assign rom_data[12556]=8'b01000000;
   assign rom_data[12557]=8'b00111100;
   assign rom_data[12558]=8'b01000000;
   assign rom_data[12559]=8'b00111101;
   assign rom_data[12560]=8'b01000000;
   assign rom_data[12561]=8'b00111110;
   assign rom_data[12562]=8'b01000000;
   assign rom_data[12563]=8'b01000000;
   assign rom_data[12564]=8'b01000000;
   assign rom_data[12565]=8'b01000001;
   assign rom_data[12566]=8'b01000000;
   assign rom_data[12567]=8'b01000010;
   assign rom_data[12568]=8'b01000000;
   assign rom_data[12569]=8'b01000100;
   assign rom_data[12570]=8'b01000000;
   assign rom_data[12571]=8'b01000101;
   assign rom_data[12572]=8'b01000000;
   assign rom_data[12573]=8'b01000110;
   assign rom_data[12574]=8'b01000000;
   assign rom_data[12575]=8'b01001000;
   assign rom_data[12576]=8'b01000000;
   assign rom_data[12577]=8'b01001001;
   assign rom_data[12578]=8'b01000000;
   assign rom_data[12579]=8'b01001010;
   assign rom_data[12580]=8'b00111111;
   assign rom_data[12581]=8'b01001100;
   assign rom_data[12582]=8'b00111111;
   assign rom_data[12583]=8'b01001101;
   assign rom_data[12584]=8'b00111111;
   assign rom_data[12585]=8'b01001110;
   assign rom_data[12586]=8'b00111111;
   assign rom_data[12587]=8'b01010000;
   assign rom_data[12588]=8'b00111111;
   assign rom_data[12589]=8'b01010001;
   assign rom_data[12590]=8'b00111111;
   assign rom_data[12591]=8'b01010011;
   assign rom_data[12592]=8'b00111111;
   assign rom_data[12593]=8'b01010100;
   assign rom_data[12594]=8'b00111111;
   assign rom_data[12595]=8'b01010101;
   assign rom_data[12596]=8'b00111111;
   assign rom_data[12597]=8'b01010111;
   assign rom_data[12598]=8'b00111111;
   assign rom_data[12599]=8'b01011000;
   assign rom_data[12600]=8'b00111111;
   assign rom_data[12601]=8'b01011010;
   assign rom_data[12602]=8'b00111111;
   assign rom_data[12603]=8'b01011011;
   assign rom_data[12604]=8'b00111111;
   assign rom_data[12605]=8'b01011100;
   assign rom_data[12606]=8'b00111111;
   assign rom_data[12607]=8'b01011110;
   assign rom_data[12608]=8'b00111111;
   assign rom_data[12609]=8'b01011111;
   assign rom_data[12610]=8'b00111111;
   assign rom_data[12611]=8'b01100001;
   assign rom_data[12612]=8'b00111111;
   assign rom_data[12613]=8'b01100010;
   assign rom_data[12614]=8'b00111111;
   assign rom_data[12615]=8'b01100011;
   assign rom_data[12616]=8'b00111111;
   assign rom_data[12617]=8'b01100101;
   assign rom_data[12618]=8'b00111111;
   assign rom_data[12619]=8'b01100110;
   assign rom_data[12620]=8'b00111111;
   assign rom_data[12621]=8'b01101000;
   assign rom_data[12622]=8'b00111111;
   assign rom_data[12623]=8'b01101001;
   assign rom_data[12624]=8'b00111111;
   assign rom_data[12625]=8'b01101010;
   assign rom_data[12626]=8'b00111111;
   assign rom_data[12627]=8'b01101100;
   assign rom_data[12628]=8'b00111111;
   assign rom_data[12629]=8'b01101101;
   assign rom_data[12630]=8'b00111111;
   assign rom_data[12631]=8'b01101110;
   assign rom_data[12632]=8'b00111111;
   assign rom_data[12633]=8'b01110000;
   assign rom_data[12634]=8'b00111111;
   assign rom_data[12635]=8'b01110001;
   assign rom_data[12636]=8'b00111111;
   assign rom_data[12637]=8'b01110010;
   assign rom_data[12638]=8'b00111111;
   assign rom_data[12639]=8'b01110100;
   assign rom_data[12640]=8'b00111111;
   assign rom_data[12641]=8'b01110101;
   assign rom_data[12642]=8'b00111111;
   assign rom_data[12643]=8'b01110110;
   assign rom_data[12644]=8'b00111111;
   assign rom_data[12645]=8'b01110111;
   assign rom_data[12646]=8'b00111111;
   assign rom_data[12647]=8'b01111001;
   assign rom_data[12648]=8'b00111111;
   assign rom_data[12649]=8'b01111010;
   assign rom_data[12650]=8'b00111111;
   assign rom_data[12651]=8'b01111011;
   assign rom_data[12652]=8'b00111111;
   assign rom_data[12653]=8'b01111100;
   assign rom_data[12654]=8'b00111111;
   assign rom_data[12655]=8'b01111101;
   assign rom_data[12656]=8'b00111111;
   assign rom_data[12657]=8'b01111110;
   assign rom_data[12658]=8'b00111111;
   assign rom_data[12659]=8'b01111111;
   assign rom_data[12660]=8'b00111111;
   assign rom_data[12661]=8'b10000000;
   assign rom_data[12662]=8'b00111110;
   assign rom_data[12663]=8'b10000001;
   assign rom_data[12664]=8'b00111110;
   assign rom_data[12665]=8'b10000010;
   assign rom_data[12666]=8'b00111110;
   assign rom_data[12667]=8'b10000011;
   assign rom_data[12668]=8'b00111110;
   assign rom_data[12669]=8'b10000100;
   assign rom_data[12670]=8'b00111110;
   assign rom_data[12671]=8'b10000101;
   assign rom_data[12672]=8'b00111110;
   assign rom_data[12673]=8'b10000110;
   assign rom_data[12674]=8'b00111110;
   assign rom_data[12675]=8'b10000110;
   assign rom_data[12676]=8'b00111110;
   assign rom_data[12677]=8'b10000111;
   assign rom_data[12678]=8'b00111110;
   assign rom_data[12679]=8'b10001000;
   assign rom_data[12680]=8'b00111110;
   assign rom_data[12681]=8'b10001000;
   assign rom_data[12682]=8'b00111110;
   assign rom_data[12683]=8'b10001001;
   assign rom_data[12684]=8'b00111110;
   assign rom_data[12685]=8'b10001001;
   assign rom_data[12686]=8'b00111110;
   assign rom_data[12687]=8'b10001001;
   assign rom_data[12688]=8'b00111110;
   assign rom_data[12689]=8'b10001010;
   assign rom_data[12690]=8'b00111110;
   assign rom_data[12691]=8'b10001010;
   assign rom_data[12692]=8'b00111110;
   assign rom_data[12693]=8'b10001010;
   assign rom_data[12694]=8'b00111110;
   assign rom_data[12695]=8'b10001010;
   assign rom_data[12696]=8'b00111110;
   assign rom_data[12697]=8'b10001010;
   assign rom_data[12698]=8'b00111110;
   assign rom_data[12699]=8'b10001001;
   assign rom_data[12700]=8'b00111110;
   assign rom_data[12701]=8'b10001001;
   assign rom_data[12702]=8'b00111110;
   assign rom_data[12703]=8'b10001001;
   assign rom_data[12704]=8'b00111110;
   assign rom_data[12705]=8'b10001000;
   assign rom_data[12706]=8'b00111110;
   assign rom_data[12707]=8'b10001000;
   assign rom_data[12708]=8'b00111110;
   assign rom_data[12709]=8'b10000111;
   assign rom_data[12710]=8'b00111110;
   assign rom_data[12711]=8'b10000111;
   assign rom_data[12712]=8'b00111110;
   assign rom_data[12713]=8'b10000110;
   assign rom_data[12714]=8'b00111110;
   assign rom_data[12715]=8'b10000101;
   assign rom_data[12716]=8'b00111110;
   assign rom_data[12717]=8'b10000100;
   assign rom_data[12718]=8'b00111110;
   assign rom_data[12719]=8'b10000011;
   assign rom_data[12720]=8'b00111110;
   assign rom_data[12721]=8'b10000011;
   assign rom_data[12722]=8'b00111110;
   assign rom_data[12723]=8'b10000010;
   assign rom_data[12724]=8'b00111110;
   assign rom_data[12725]=8'b10000001;
   assign rom_data[12726]=8'b00111110;
   assign rom_data[12727]=8'b01111111;
   assign rom_data[12728]=8'b00111101;
   assign rom_data[12729]=8'b01111110;
   assign rom_data[12730]=8'b00111101;
   assign rom_data[12731]=8'b01111101;
   assign rom_data[12732]=8'b00111101;
   assign rom_data[12733]=8'b01111100;
   assign rom_data[12734]=8'b00111101;
   assign rom_data[12735]=8'b01111011;
   assign rom_data[12736]=8'b00111101;
   assign rom_data[12737]=8'b01111010;
   assign rom_data[12738]=8'b00111101;
   assign rom_data[12739]=8'b01111001;
   assign rom_data[12740]=8'b00111101;
   assign rom_data[12741]=8'b01110111;
   assign rom_data[12742]=8'b00111101;
   assign rom_data[12743]=8'b01110110;
   assign rom_data[12744]=8'b00111101;
   assign rom_data[12745]=8'b01110101;
   assign rom_data[12746]=8'b00111101;
   assign rom_data[12747]=8'b01110100;
   assign rom_data[12748]=8'b00111101;
   assign rom_data[12749]=8'b01110010;
   assign rom_data[12750]=8'b00111101;
   assign rom_data[12751]=8'b01110001;
   assign rom_data[12752]=8'b00111101;
   assign rom_data[12753]=8'b01110000;
   assign rom_data[12754]=8'b00111101;
   assign rom_data[12755]=8'b01101110;
   assign rom_data[12756]=8'b00111101;
   assign rom_data[12757]=8'b01101101;
   assign rom_data[12758]=8'b00111101;
   assign rom_data[12759]=8'b01101100;
   assign rom_data[12760]=8'b00111101;
   assign rom_data[12761]=8'b01101010;
   assign rom_data[12762]=8'b00111101;
   assign rom_data[12763]=8'b01101001;
   assign rom_data[12764]=8'b00111101;
   assign rom_data[12765]=8'b01100111;
   assign rom_data[12766]=8'b00111101;
   assign rom_data[12767]=8'b01100110;
   assign rom_data[12768]=8'b00111101;
   assign rom_data[12769]=8'b01100101;
   assign rom_data[12770]=8'b00111101;
   assign rom_data[12771]=8'b01100011;
   assign rom_data[12772]=8'b00111101;
   assign rom_data[12773]=8'b01100010;
   assign rom_data[12774]=8'b00111101;
   assign rom_data[12775]=8'b01100000;
   assign rom_data[12776]=8'b00111101;
   assign rom_data[12777]=8'b01011111;
   assign rom_data[12778]=8'b00111101;
   assign rom_data[12779]=8'b01011110;
   assign rom_data[12780]=8'b00111101;
   assign rom_data[12781]=8'b01011100;
   assign rom_data[12782]=8'b00111101;
   assign rom_data[12783]=8'b01011011;
   assign rom_data[12784]=8'b00111101;
   assign rom_data[12785]=8'b01011001;
   assign rom_data[12786]=8'b00111101;
   assign rom_data[12787]=8'b01011000;
   assign rom_data[12788]=8'b00111101;
   assign rom_data[12789]=8'b01010111;
   assign rom_data[12790]=8'b00111101;
   assign rom_data[12791]=8'b01010101;
   assign rom_data[12792]=8'b00111101;
   assign rom_data[12793]=8'b01010100;
   assign rom_data[12794]=8'b00111101;
   assign rom_data[12795]=8'b01010010;
   assign rom_data[12796]=8'b00111101;
   assign rom_data[12797]=8'b01010001;
   assign rom_data[12798]=8'b00111101;
   assign rom_data[12799]=8'b01010000;
   assign rom_data[12800]=8'b00111101;
   assign rom_data[12801]=8'b01001110;
   assign rom_data[12802]=8'b00111101;
   assign rom_data[12803]=8'b01001101;
   assign rom_data[12804]=8'b00111101;
   assign rom_data[12805]=8'b01001100;
   assign rom_data[12806]=8'b00111101;
   assign rom_data[12807]=8'b01001010;
   assign rom_data[12808]=8'b00111101;
   assign rom_data[12809]=8'b01001001;
   assign rom_data[12810]=8'b00111101;
   assign rom_data[12811]=8'b01000111;
   assign rom_data[12812]=8'b00111100;
   assign rom_data[12813]=8'b01000110;
   assign rom_data[12814]=8'b00111100;
   assign rom_data[12815]=8'b01000101;
   assign rom_data[12816]=8'b00111100;
   assign rom_data[12817]=8'b01000100;
   assign rom_data[12818]=8'b00111100;
   assign rom_data[12819]=8'b01000010;
   assign rom_data[12820]=8'b00111100;
   assign rom_data[12821]=8'b01000001;
   assign rom_data[12822]=8'b00111100;
   assign rom_data[12823]=8'b01000000;
   assign rom_data[12824]=8'b00111100;
   assign rom_data[12825]=8'b00111110;
   assign rom_data[12826]=8'b00111100;
   assign rom_data[12827]=8'b00111101;
   assign rom_data[12828]=8'b00111100;
   assign rom_data[12829]=8'b00111100;
   assign rom_data[12830]=8'b00111100;
   assign rom_data[12831]=8'b00111011;
   assign rom_data[12832]=8'b00111100;
   assign rom_data[12833]=8'b00111010;
   assign rom_data[12834]=8'b00111100;
   assign rom_data[12835]=8'b00111001;
   assign rom_data[12836]=8'b00111100;
   assign rom_data[12837]=8'b00110111;
   assign rom_data[12838]=8'b00111100;
   assign rom_data[12839]=8'b00110110;
   assign rom_data[12840]=8'b00111100;
   assign rom_data[12841]=8'b00110101;
   assign rom_data[12842]=8'b00111100;
   assign rom_data[12843]=8'b00110100;
   assign rom_data[12844]=8'b00111100;
   assign rom_data[12845]=8'b00110011;
   assign rom_data[12846]=8'b00111100;
   assign rom_data[12847]=8'b00110011;
   assign rom_data[12848]=8'b00111100;
   assign rom_data[12849]=8'b00110010;
   assign rom_data[12850]=8'b00111100;
   assign rom_data[12851]=8'b00110001;
   assign rom_data[12852]=8'b00111100;
   assign rom_data[12853]=8'b00110000;
   assign rom_data[12854]=8'b00111100;
   assign rom_data[12855]=8'b00101111;
   assign rom_data[12856]=8'b00111100;
   assign rom_data[12857]=8'b00101111;
   assign rom_data[12858]=8'b00111100;
   assign rom_data[12859]=8'b00101110;
   assign rom_data[12860]=8'b00111100;
   assign rom_data[12861]=8'b00101110;
   assign rom_data[12862]=8'b00111100;
   assign rom_data[12863]=8'b00101101;
   assign rom_data[12864]=8'b00111100;
   assign rom_data[12865]=8'b00101101;
   assign rom_data[12866]=8'b00111100;
   assign rom_data[12867]=8'b00101100;
   assign rom_data[12868]=8'b00111100;
   assign rom_data[12869]=8'b00101100;
   assign rom_data[12870]=8'b00111100;
   assign rom_data[12871]=8'b00101100;
   assign rom_data[12872]=8'b00111100;
   assign rom_data[12873]=8'b00101100;
   assign rom_data[12874]=8'b00111100;
   assign rom_data[12875]=8'b00101100;
   assign rom_data[12876]=8'b00111100;
   assign rom_data[12877]=8'b00101100;
   assign rom_data[12878]=8'b00111100;
   assign rom_data[12879]=8'b00101100;
   assign rom_data[12880]=8'b00111011;
   assign rom_data[12881]=8'b00101101;
   assign rom_data[12882]=8'b00111011;
   assign rom_data[12883]=8'b00101101;
   assign rom_data[12884]=8'b00111011;
   assign rom_data[12885]=8'b00101101;
   assign rom_data[12886]=8'b00111011;
   assign rom_data[12887]=8'b00101110;
   assign rom_data[12888]=8'b00111011;
   assign rom_data[12889]=8'b00101111;
   assign rom_data[12890]=8'b00111011;
   assign rom_data[12891]=8'b00101111;
   assign rom_data[12892]=8'b00111011;
   assign rom_data[12893]=8'b00110000;
   assign rom_data[12894]=8'b00111011;
   assign rom_data[12895]=8'b00110001;
   assign rom_data[12896]=8'b00111011;
   assign rom_data[12897]=8'b00110010;
   assign rom_data[12898]=8'b00111011;
   assign rom_data[12899]=8'b00110010;
   assign rom_data[12900]=8'b00111011;
   assign rom_data[12901]=8'b00110011;
   assign rom_data[12902]=8'b00111011;
   assign rom_data[12903]=8'b00110100;
   assign rom_data[12904]=8'b00111011;
   assign rom_data[12905]=8'b00110101;
   assign rom_data[12906]=8'b00111011;
   assign rom_data[12907]=8'b00110110;
   assign rom_data[12908]=8'b00111011;
   assign rom_data[12909]=8'b00110111;
   assign rom_data[12910]=8'b00111011;
   assign rom_data[12911]=8'b00111001;
   assign rom_data[12912]=8'b00111011;
   assign rom_data[12913]=8'b00111010;
   assign rom_data[12914]=8'b00111011;
   assign rom_data[12915]=8'b00111011;
   assign rom_data[12916]=8'b00111011;
   assign rom_data[12917]=8'b00111100;
   assign rom_data[12918]=8'b00111011;
   assign rom_data[12919]=8'b00111101;
   assign rom_data[12920]=8'b00111011;
   assign rom_data[12921]=8'b00111110;
   assign rom_data[12922]=8'b00111011;
   assign rom_data[12923]=8'b01000000;
   assign rom_data[12924]=8'b00111011;
   assign rom_data[12925]=8'b01000001;
   assign rom_data[12926]=8'b00111011;
   assign rom_data[12927]=8'b01000010;
   assign rom_data[12928]=8'b00111011;
   assign rom_data[12929]=8'b01000100;
   assign rom_data[12930]=8'b00111011;
   assign rom_data[12931]=8'b01000101;
   assign rom_data[12932]=8'b00111011;
   assign rom_data[12933]=8'b01000110;
   assign rom_data[12934]=8'b00111011;
   assign rom_data[12935]=8'b01001000;
   assign rom_data[12936]=8'b00111011;
   assign rom_data[12937]=8'b01001001;
   assign rom_data[12938]=8'b00111011;
   assign rom_data[12939]=8'b01001010;
   assign rom_data[12940]=8'b00111011;
   assign rom_data[12941]=8'b01001100;
   assign rom_data[12942]=8'b00111011;
   assign rom_data[12943]=8'b01001101;
   assign rom_data[12944]=8'b00111011;
   assign rom_data[12945]=8'b01001110;
   assign rom_data[12946]=8'b00111011;
   assign rom_data[12947]=8'b01010000;
   assign rom_data[12948]=8'b00111011;
   assign rom_data[12949]=8'b01010001;
   assign rom_data[12950]=8'b00111011;
   assign rom_data[12951]=8'b01010011;
   assign rom_data[12952]=8'b00111011;
   assign rom_data[12953]=8'b01010100;
   assign rom_data[12954]=8'b00111011;
   assign rom_data[12955]=8'b01010101;
   assign rom_data[12956]=8'b00111011;
   assign rom_data[12957]=8'b01010111;
   assign rom_data[12958]=8'b00111010;
   assign rom_data[12959]=8'b01011000;
   assign rom_data[12960]=8'b00111010;
   assign rom_data[12961]=8'b01011010;
   assign rom_data[12962]=8'b00111010;
   assign rom_data[12963]=8'b01011011;
   assign rom_data[12964]=8'b00111010;
   assign rom_data[12965]=8'b01011100;
   assign rom_data[12966]=8'b00111010;
   assign rom_data[12967]=8'b01011110;
   assign rom_data[12968]=8'b00111010;
   assign rom_data[12969]=8'b01011111;
   assign rom_data[12970]=8'b00111010;
   assign rom_data[12971]=8'b01100001;
   assign rom_data[12972]=8'b00111010;
   assign rom_data[12973]=8'b01100010;
   assign rom_data[12974]=8'b00111010;
   assign rom_data[12975]=8'b01100011;
   assign rom_data[12976]=8'b00111010;
   assign rom_data[12977]=8'b01100101;
   assign rom_data[12978]=8'b00111010;
   assign rom_data[12979]=8'b01100110;
   assign rom_data[12980]=8'b00111010;
   assign rom_data[12981]=8'b01101000;
   assign rom_data[12982]=8'b00111010;
   assign rom_data[12983]=8'b01101001;
   assign rom_data[12984]=8'b00111010;
   assign rom_data[12985]=8'b01101010;
   assign rom_data[12986]=8'b00111010;
   assign rom_data[12987]=8'b01101100;
   assign rom_data[12988]=8'b00111010;
   assign rom_data[12989]=8'b01101101;
   assign rom_data[12990]=8'b00111010;
   assign rom_data[12991]=8'b01101110;
   assign rom_data[12992]=8'b00111010;
   assign rom_data[12993]=8'b01110000;
   assign rom_data[12994]=8'b00111010;
   assign rom_data[12995]=8'b01110001;
   assign rom_data[12996]=8'b00111010;
   assign rom_data[12997]=8'b01110010;
   assign rom_data[12998]=8'b00111010;
   assign rom_data[12999]=8'b01110100;
   assign rom_data[13000]=8'b00111010;
   assign rom_data[13001]=8'b01110101;
   assign rom_data[13002]=8'b00111010;
   assign rom_data[13003]=8'b01110110;
   assign rom_data[13004]=8'b00111010;
   assign rom_data[13005]=8'b01110111;
   assign rom_data[13006]=8'b00111010;
   assign rom_data[13007]=8'b01111001;
   assign rom_data[13008]=8'b00111010;
   assign rom_data[13009]=8'b01111010;
   assign rom_data[13010]=8'b00111010;
   assign rom_data[13011]=8'b01111011;
   assign rom_data[13012]=8'b00111010;
   assign rom_data[13013]=8'b01111100;
   assign rom_data[13014]=8'b00111010;
   assign rom_data[13015]=8'b01111101;
   assign rom_data[13016]=8'b00111010;
   assign rom_data[13017]=8'b01111110;
   assign rom_data[13018]=8'b00111010;
   assign rom_data[13019]=8'b01111111;
   assign rom_data[13020]=8'b00111010;
   assign rom_data[13021]=8'b10000000;
   assign rom_data[13022]=8'b00111010;
   assign rom_data[13023]=8'b10000001;
   assign rom_data[13024]=8'b00111010;
   assign rom_data[13025]=8'b10000010;
   assign rom_data[13026]=8'b00111010;
   assign rom_data[13027]=8'b10000011;
   assign rom_data[13028]=8'b00111010;
   assign rom_data[13029]=8'b10000100;
   assign rom_data[13030]=8'b00111010;
   assign rom_data[13031]=8'b10000101;
   assign rom_data[13032]=8'b00111010;
   assign rom_data[13033]=8'b10000110;
   assign rom_data[13034]=8'b00111010;
   assign rom_data[13035]=8'b10000110;
   assign rom_data[13036]=8'b00111001;
   assign rom_data[13037]=8'b10000111;
   assign rom_data[13038]=8'b00111001;
   assign rom_data[13039]=8'b10001000;
   assign rom_data[13040]=8'b00111001;
   assign rom_data[13041]=8'b10001000;
   assign rom_data[13042]=8'b00111001;
   assign rom_data[13043]=8'b10001001;
   assign rom_data[13044]=8'b00111001;
   assign rom_data[13045]=8'b10001001;
   assign rom_data[13046]=8'b00111001;
   assign rom_data[13047]=8'b10001001;
   assign rom_data[13048]=8'b00111001;
   assign rom_data[13049]=8'b10001010;
   assign rom_data[13050]=8'b00111001;
   assign rom_data[13051]=8'b10001010;
   assign rom_data[13052]=8'b00111001;
   assign rom_data[13053]=8'b10001010;
   assign rom_data[13054]=8'b00111001;
   assign rom_data[13055]=8'b10001010;
   assign rom_data[13056]=8'b00111001;
   assign rom_data[13057]=8'b10001010;
   assign rom_data[13058]=8'b00111001;
   assign rom_data[13059]=8'b10001001;
   assign rom_data[13060]=8'b00111001;
   assign rom_data[13061]=8'b10001001;
   assign rom_data[13062]=8'b00111001;
   assign rom_data[13063]=8'b10001001;
   assign rom_data[13064]=8'b00111001;
   assign rom_data[13065]=8'b10001000;
   assign rom_data[13066]=8'b00111001;
   assign rom_data[13067]=8'b10001000;
   assign rom_data[13068]=8'b00111001;
   assign rom_data[13069]=8'b10000111;
   assign rom_data[13070]=8'b00111001;
   assign rom_data[13071]=8'b10000111;
   assign rom_data[13072]=8'b00111001;
   assign rom_data[13073]=8'b10000110;
   assign rom_data[13074]=8'b00111001;
   assign rom_data[13075]=8'b10000101;
   assign rom_data[13076]=8'b00111001;
   assign rom_data[13077]=8'b10000100;
   assign rom_data[13078]=8'b00111001;
   assign rom_data[13079]=8'b10000011;
   assign rom_data[13080]=8'b00111001;
   assign rom_data[13081]=8'b10000011;
   assign rom_data[13082]=8'b00111001;
   assign rom_data[13083]=8'b10000010;
   assign rom_data[13084]=8'b00111001;
   assign rom_data[13085]=8'b10000001;
   assign rom_data[13086]=8'b00111001;
   assign rom_data[13087]=8'b01111111;
   assign rom_data[13088]=8'b00111001;
   assign rom_data[13089]=8'b01111110;
   assign rom_data[13090]=8'b00111001;
   assign rom_data[13091]=8'b01111101;
   assign rom_data[13092]=8'b00111001;
   assign rom_data[13093]=8'b01111100;
   assign rom_data[13094]=8'b00111001;
   assign rom_data[13095]=8'b01111011;
   assign rom_data[13096]=8'b00111001;
   assign rom_data[13097]=8'b01111010;
   assign rom_data[13098]=8'b00111001;
   assign rom_data[13099]=8'b01111001;
   assign rom_data[13100]=8'b00111001;
   assign rom_data[13101]=8'b01110111;
   assign rom_data[13102]=8'b00111001;
   assign rom_data[13103]=8'b01110110;
   assign rom_data[13104]=8'b00111000;
   assign rom_data[13105]=8'b01110101;
   assign rom_data[13106]=8'b00111000;
   assign rom_data[13107]=8'b01110100;
   assign rom_data[13108]=8'b00111000;
   assign rom_data[13109]=8'b01110010;
   assign rom_data[13110]=8'b00111000;
   assign rom_data[13111]=8'b01110001;
   assign rom_data[13112]=8'b00111000;
   assign rom_data[13113]=8'b01110000;
   assign rom_data[13114]=8'b00111000;
   assign rom_data[13115]=8'b01101110;
   assign rom_data[13116]=8'b00111000;
   assign rom_data[13117]=8'b01101101;
   assign rom_data[13118]=8'b00111000;
   assign rom_data[13119]=8'b01101100;
   assign rom_data[13120]=8'b00111000;
   assign rom_data[13121]=8'b01101010;
   assign rom_data[13122]=8'b00111000;
   assign rom_data[13123]=8'b01101001;
   assign rom_data[13124]=8'b00111000;
   assign rom_data[13125]=8'b01100111;
   assign rom_data[13126]=8'b00111000;
   assign rom_data[13127]=8'b01100110;
   assign rom_data[13128]=8'b00111000;
   assign rom_data[13129]=8'b01100101;
   assign rom_data[13130]=8'b00111000;
   assign rom_data[13131]=8'b01100011;
   assign rom_data[13132]=8'b00111000;
   assign rom_data[13133]=8'b01100010;
   assign rom_data[13134]=8'b00111000;
   assign rom_data[13135]=8'b01100000;
   assign rom_data[13136]=8'b00111000;
   assign rom_data[13137]=8'b01011111;
   assign rom_data[13138]=8'b00111000;
   assign rom_data[13139]=8'b01011110;
   assign rom_data[13140]=8'b00111000;
   assign rom_data[13141]=8'b01011100;
   assign rom_data[13142]=8'b00111000;
   assign rom_data[13143]=8'b01011011;
   assign rom_data[13144]=8'b00111000;
   assign rom_data[13145]=8'b01011001;
   assign rom_data[13146]=8'b00111000;
   assign rom_data[13147]=8'b01011000;
   assign rom_data[13148]=8'b00111000;
   assign rom_data[13149]=8'b01010111;
   assign rom_data[13150]=8'b00111000;
   assign rom_data[13151]=8'b01010101;
   assign rom_data[13152]=8'b00111000;
   assign rom_data[13153]=8'b01010100;
   assign rom_data[13154]=8'b00111000;
   assign rom_data[13155]=8'b01010010;
   assign rom_data[13156]=8'b00111000;
   assign rom_data[13157]=8'b01010001;
   assign rom_data[13158]=8'b00111000;
   assign rom_data[13159]=8'b01010000;
   assign rom_data[13160]=8'b00111000;
   assign rom_data[13161]=8'b01001110;
   assign rom_data[13162]=8'b00111000;
   assign rom_data[13163]=8'b01001101;
   assign rom_data[13164]=8'b00111000;
   assign rom_data[13165]=8'b01001100;
   assign rom_data[13166]=8'b00111000;
   assign rom_data[13167]=8'b01001010;
   assign rom_data[13168]=8'b00111000;
   assign rom_data[13169]=8'b01001001;
   assign rom_data[13170]=8'b00111000;
   assign rom_data[13171]=8'b01000111;
   assign rom_data[13172]=8'b00111000;
   assign rom_data[13173]=8'b01000110;
   assign rom_data[13174]=8'b00111000;
   assign rom_data[13175]=8'b01000101;
   assign rom_data[13176]=8'b00111000;
   assign rom_data[13177]=8'b01000100;
   assign rom_data[13178]=8'b00111000;
   assign rom_data[13179]=8'b01000010;
   assign rom_data[13180]=8'b00111000;
   assign rom_data[13181]=8'b01000001;
   assign rom_data[13182]=8'b00111000;
   assign rom_data[13183]=8'b01000000;
   assign rom_data[13184]=8'b00111000;
   assign rom_data[13185]=8'b00111110;
   assign rom_data[13186]=8'b00111000;
   assign rom_data[13187]=8'b00111101;
   assign rom_data[13188]=8'b00110111;
   assign rom_data[13189]=8'b00111100;
   assign rom_data[13190]=8'b00110111;
   assign rom_data[13191]=8'b00111011;
   assign rom_data[13192]=8'b00110111;
   assign rom_data[13193]=8'b00111010;
   assign rom_data[13194]=8'b00110111;
   assign rom_data[13195]=8'b00111001;
   assign rom_data[13196]=8'b00110111;
   assign rom_data[13197]=8'b00110111;
   assign rom_data[13198]=8'b00110111;
   assign rom_data[13199]=8'b00110110;
   assign rom_data[13200]=8'b00110111;
   assign rom_data[13201]=8'b00110101;
   assign rom_data[13202]=8'b00110111;
   assign rom_data[13203]=8'b00110100;
   assign rom_data[13204]=8'b00110111;
   assign rom_data[13205]=8'b00110011;
   assign rom_data[13206]=8'b00110111;
   assign rom_data[13207]=8'b00110011;
   assign rom_data[13208]=8'b00110111;
   assign rom_data[13209]=8'b00110010;
   assign rom_data[13210]=8'b00110111;
   assign rom_data[13211]=8'b00110001;
   assign rom_data[13212]=8'b00110111;
   assign rom_data[13213]=8'b00110000;
   assign rom_data[13214]=8'b00110111;
   assign rom_data[13215]=8'b00101111;
   assign rom_data[13216]=8'b00110111;
   assign rom_data[13217]=8'b00101111;
   assign rom_data[13218]=8'b00110111;
   assign rom_data[13219]=8'b00101110;
   assign rom_data[13220]=8'b00110111;
   assign rom_data[13221]=8'b00101110;
   assign rom_data[13222]=8'b00110111;
   assign rom_data[13223]=8'b00101101;
   assign rom_data[13224]=8'b00110111;
   assign rom_data[13225]=8'b00101101;
   assign rom_data[13226]=8'b00110111;
   assign rom_data[13227]=8'b00101100;
   assign rom_data[13228]=8'b00110111;
   assign rom_data[13229]=8'b00101100;
   assign rom_data[13230]=8'b00110111;
   assign rom_data[13231]=8'b00101100;
   assign rom_data[13232]=8'b00110111;
   assign rom_data[13233]=8'b00101100;
   assign rom_data[13234]=8'b00110111;
   assign rom_data[13235]=8'b00101100;
   assign rom_data[13236]=8'b00110111;
   assign rom_data[13237]=8'b00101100;
   assign rom_data[13238]=8'b00110111;
   assign rom_data[13239]=8'b00101100;
   assign rom_data[13240]=8'b00110111;
   assign rom_data[13241]=8'b00101101;
   assign rom_data[13242]=8'b00110111;
   assign rom_data[13243]=8'b00101101;
   assign rom_data[13244]=8'b00110111;
   assign rom_data[13245]=8'b00101101;
   assign rom_data[13246]=8'b00110111;
   assign rom_data[13247]=8'b00101110;
   assign rom_data[13248]=8'b00110111;
   assign rom_data[13249]=8'b00101111;
   assign rom_data[13250]=8'b00110111;
   assign rom_data[13251]=8'b00101111;
   assign rom_data[13252]=8'b00110111;
   assign rom_data[13253]=8'b00110000;
   assign rom_data[13254]=8'b00110110;
   assign rom_data[13255]=8'b00110001;
   assign rom_data[13256]=8'b00110110;
   assign rom_data[13257]=8'b00110010;
   assign rom_data[13258]=8'b00110110;
   assign rom_data[13259]=8'b00110010;
   assign rom_data[13260]=8'b00110110;
   assign rom_data[13261]=8'b00110011;
   assign rom_data[13262]=8'b00110110;
   assign rom_data[13263]=8'b00110100;
   assign rom_data[13264]=8'b00110110;
   assign rom_data[13265]=8'b00110101;
   assign rom_data[13266]=8'b00110110;
   assign rom_data[13267]=8'b00110110;
   assign rom_data[13268]=8'b00110110;
   assign rom_data[13269]=8'b00110111;
   assign rom_data[13270]=8'b00110110;
   assign rom_data[13271]=8'b00111001;
   assign rom_data[13272]=8'b00110110;
   assign rom_data[13273]=8'b00111010;
   assign rom_data[13274]=8'b00110110;
   assign rom_data[13275]=8'b00111011;
   assign rom_data[13276]=8'b00110110;
   assign rom_data[13277]=8'b00111100;
   assign rom_data[13278]=8'b00110110;
   assign rom_data[13279]=8'b00111101;
   assign rom_data[13280]=8'b00110110;
   assign rom_data[13281]=8'b00111110;
   assign rom_data[13282]=8'b00110110;
   assign rom_data[13283]=8'b01000000;
   assign rom_data[13284]=8'b00110110;
   assign rom_data[13285]=8'b01000001;
   assign rom_data[13286]=8'b00110110;
   assign rom_data[13287]=8'b01000010;
   assign rom_data[13288]=8'b00110110;
   assign rom_data[13289]=8'b01000100;
   assign rom_data[13290]=8'b00110110;
   assign rom_data[13291]=8'b01000101;
   assign rom_data[13292]=8'b00110110;
   assign rom_data[13293]=8'b01000110;
   assign rom_data[13294]=8'b00110110;
   assign rom_data[13295]=8'b01001000;
   assign rom_data[13296]=8'b00110110;
   assign rom_data[13297]=8'b01001001;
   assign rom_data[13298]=8'b00110110;
   assign rom_data[13299]=8'b01001010;
   assign rom_data[13300]=8'b00110110;
   assign rom_data[13301]=8'b01001100;
   assign rom_data[13302]=8'b00110110;
   assign rom_data[13303]=8'b01001101;
   assign rom_data[13304]=8'b00110110;
   assign rom_data[13305]=8'b01001110;
   assign rom_data[13306]=8'b00110110;
   assign rom_data[13307]=8'b01010000;
   assign rom_data[13308]=8'b00110110;
   assign rom_data[13309]=8'b01010001;
   assign rom_data[13310]=8'b00110110;
   assign rom_data[13311]=8'b01010011;
   assign rom_data[13312]=8'b00110110;
   assign rom_data[13313]=8'b01010100;
   assign rom_data[13314]=8'b00110110;
   assign rom_data[13315]=8'b01010101;
   assign rom_data[13316]=8'b00110110;
   assign rom_data[13317]=8'b01010111;
   assign rom_data[13318]=8'b00110110;
   assign rom_data[13319]=8'b01011000;
   assign rom_data[13320]=8'b00110110;
   assign rom_data[13321]=8'b01011010;
   assign rom_data[13322]=8'b00110110;
   assign rom_data[13323]=8'b01011011;
   assign rom_data[13324]=8'b00110110;
   assign rom_data[13325]=8'b01011100;
   assign rom_data[13326]=8'b00110110;
   assign rom_data[13327]=8'b01011110;
   assign rom_data[13328]=8'b00110110;
   assign rom_data[13329]=8'b01011111;
   assign rom_data[13330]=8'b00110110;
   assign rom_data[13331]=8'b01100001;
   assign rom_data[13332]=8'b00110110;
   assign rom_data[13333]=8'b01100010;
   assign rom_data[13334]=8'b00110101;
   assign rom_data[13335]=8'b01100011;
   assign rom_data[13336]=8'b00110101;
   assign rom_data[13337]=8'b01100101;
   assign rom_data[13338]=8'b00110101;
   assign rom_data[13339]=8'b01100110;
   assign rom_data[13340]=8'b00110101;
   assign rom_data[13341]=8'b01101000;
   assign rom_data[13342]=8'b00110101;
   assign rom_data[13343]=8'b01101001;
   assign rom_data[13344]=8'b00110101;
   assign rom_data[13345]=8'b01101010;
   assign rom_data[13346]=8'b00110101;
   assign rom_data[13347]=8'b01101100;
   assign rom_data[13348]=8'b00110101;
   assign rom_data[13349]=8'b01101101;
   assign rom_data[13350]=8'b00110101;
   assign rom_data[13351]=8'b01101110;
   assign rom_data[13352]=8'b00110101;
   assign rom_data[13353]=8'b01110000;
   assign rom_data[13354]=8'b00110101;
   assign rom_data[13355]=8'b01110001;
   assign rom_data[13356]=8'b00110101;
   assign rom_data[13357]=8'b01110010;
   assign rom_data[13358]=8'b00110101;
   assign rom_data[13359]=8'b01110100;
   assign rom_data[13360]=8'b00110101;
   assign rom_data[13361]=8'b01110101;
   assign rom_data[13362]=8'b00110101;
   assign rom_data[13363]=8'b01110110;
   assign rom_data[13364]=8'b00110101;
   assign rom_data[13365]=8'b01110111;
   assign rom_data[13366]=8'b00110101;
   assign rom_data[13367]=8'b01111001;
   assign rom_data[13368]=8'b00110101;
   assign rom_data[13369]=8'b01111010;
   assign rom_data[13370]=8'b00110101;
   assign rom_data[13371]=8'b01111011;
   assign rom_data[13372]=8'b00110101;
   assign rom_data[13373]=8'b01111100;
   assign rom_data[13374]=8'b00110101;
   assign rom_data[13375]=8'b01111101;
   assign rom_data[13376]=8'b00110101;
   assign rom_data[13377]=8'b01111110;
   assign rom_data[13378]=8'b00110101;
   assign rom_data[13379]=8'b01111111;
   assign rom_data[13380]=8'b00110101;
   assign rom_data[13381]=8'b10000000;
   assign rom_data[13382]=8'b00110101;
   assign rom_data[13383]=8'b10000001;
   assign rom_data[13384]=8'b00110101;
   assign rom_data[13385]=8'b10000010;
   assign rom_data[13386]=8'b00110101;
   assign rom_data[13387]=8'b10000011;
   assign rom_data[13388]=8'b00110101;
   assign rom_data[13389]=8'b10000100;
   assign rom_data[13390]=8'b00110101;
   assign rom_data[13391]=8'b10000101;
   assign rom_data[13392]=8'b00110101;
   assign rom_data[13393]=8'b10000110;
   assign rom_data[13394]=8'b00110101;
   assign rom_data[13395]=8'b10000110;
   assign rom_data[13396]=8'b00110101;
   assign rom_data[13397]=8'b10000111;
   assign rom_data[13398]=8'b00110101;
   assign rom_data[13399]=8'b10001000;
   assign rom_data[13400]=8'b00110101;
   assign rom_data[13401]=8'b10001000;
   assign rom_data[13402]=8'b00110101;
   assign rom_data[13403]=8'b10001001;
   assign rom_data[13404]=8'b00110101;
   assign rom_data[13405]=8'b10001001;
   assign rom_data[13406]=8'b00110101;
   assign rom_data[13407]=8'b10001001;
   assign rom_data[13408]=8'b00110100;
   assign rom_data[13409]=8'b10001010;
   assign rom_data[13410]=8'b00110100;
   assign rom_data[13411]=8'b10001010;
   assign rom_data[13412]=8'b00110100;
   assign rom_data[13413]=8'b10001010;
   assign rom_data[13414]=8'b00110100;
   assign rom_data[13415]=8'b10001010;
   assign rom_data[13416]=8'b00110100;
   assign rom_data[13417]=8'b10001010;
   assign rom_data[13418]=8'b00110100;
   assign rom_data[13419]=8'b10001001;
   assign rom_data[13420]=8'b00110100;
   assign rom_data[13421]=8'b10001001;
   assign rom_data[13422]=8'b00110100;
   assign rom_data[13423]=8'b10001001;
   assign rom_data[13424]=8'b00110100;
   assign rom_data[13425]=8'b10001000;
   assign rom_data[13426]=8'b00110100;
   assign rom_data[13427]=8'b10001000;
   assign rom_data[13428]=8'b00110100;
   assign rom_data[13429]=8'b10000111;
   assign rom_data[13430]=8'b00110100;
   assign rom_data[13431]=8'b10000111;
   assign rom_data[13432]=8'b00110100;
   assign rom_data[13433]=8'b10000110;
   assign rom_data[13434]=8'b00110100;
   assign rom_data[13435]=8'b10000101;
   assign rom_data[13436]=8'b00110100;
   assign rom_data[13437]=8'b10000100;
   assign rom_data[13438]=8'b00110100;
   assign rom_data[13439]=8'b10000011;
   assign rom_data[13440]=8'b00110100;
   assign rom_data[13441]=8'b10000011;
   assign rom_data[13442]=8'b00110100;
   assign rom_data[13443]=8'b10000010;
   assign rom_data[13444]=8'b00110100;
   assign rom_data[13445]=8'b10000001;
   assign rom_data[13446]=8'b00110100;
   assign rom_data[13447]=8'b01111111;
   assign rom_data[13448]=8'b00110100;
   assign rom_data[13449]=8'b01111110;
   assign rom_data[13450]=8'b00110100;
   assign rom_data[13451]=8'b01111101;
   assign rom_data[13452]=8'b00110100;
   assign rom_data[13453]=8'b01111100;
   assign rom_data[13454]=8'b00110100;
   assign rom_data[13455]=8'b01111011;
   assign rom_data[13456]=8'b00110100;
   assign rom_data[13457]=8'b01111010;
   assign rom_data[13458]=8'b00110100;
   assign rom_data[13459]=8'b01111001;
   assign rom_data[13460]=8'b00110100;
   assign rom_data[13461]=8'b01110111;
   assign rom_data[13462]=8'b00110100;
   assign rom_data[13463]=8'b01110110;
   assign rom_data[13464]=8'b00110100;
   assign rom_data[13465]=8'b01110101;
   assign rom_data[13466]=8'b00110100;
   assign rom_data[13467]=8'b01110100;
   assign rom_data[13468]=8'b00110100;
   assign rom_data[13469]=8'b01110010;
   assign rom_data[13470]=8'b00110100;
   assign rom_data[13471]=8'b01110001;
   assign rom_data[13472]=8'b00110100;
   assign rom_data[13473]=8'b01110000;
   assign rom_data[13474]=8'b00110100;
   assign rom_data[13475]=8'b01101110;
   assign rom_data[13476]=8'b00110100;
   assign rom_data[13477]=8'b01101101;
   assign rom_data[13478]=8'b00110100;
   assign rom_data[13479]=8'b01101100;
   assign rom_data[13480]=8'b00110011;
   assign rom_data[13481]=8'b01101010;
   assign rom_data[13482]=8'b00110011;
   assign rom_data[13483]=8'b01101001;
   assign rom_data[13484]=8'b00110011;
   assign rom_data[13485]=8'b01100111;
   assign rom_data[13486]=8'b00110011;
   assign rom_data[13487]=8'b01100110;
   assign rom_data[13488]=8'b00110011;
   assign rom_data[13489]=8'b01100101;
   assign rom_data[13490]=8'b00110011;
   assign rom_data[13491]=8'b01100011;
   assign rom_data[13492]=8'b00110011;
   assign rom_data[13493]=8'b01100010;
   assign rom_data[13494]=8'b00110011;
   assign rom_data[13495]=8'b01100000;
   assign rom_data[13496]=8'b00110011;
   assign rom_data[13497]=8'b01011111;
   assign rom_data[13498]=8'b00110011;
   assign rom_data[13499]=8'b01011110;
   assign rom_data[13500]=8'b00110011;
   assign rom_data[13501]=8'b01011100;
   assign rom_data[13502]=8'b00110011;
   assign rom_data[13503]=8'b01011011;
   assign rom_data[13504]=8'b00110011;
   assign rom_data[13505]=8'b01011001;
   assign rom_data[13506]=8'b00110011;
   assign rom_data[13507]=8'b01011000;
   assign rom_data[13508]=8'b00110011;
   assign rom_data[13509]=8'b01010111;
   assign rom_data[13510]=8'b00110011;
   assign rom_data[13511]=8'b01010101;
   assign rom_data[13512]=8'b00110011;
   assign rom_data[13513]=8'b01010100;
   assign rom_data[13514]=8'b00110011;
   assign rom_data[13515]=8'b01010010;
   assign rom_data[13516]=8'b00110011;
   assign rom_data[13517]=8'b01010001;
   assign rom_data[13518]=8'b00110011;
   assign rom_data[13519]=8'b01010000;
   assign rom_data[13520]=8'b00110011;
   assign rom_data[13521]=8'b01001110;
   assign rom_data[13522]=8'b00110011;
   assign rom_data[13523]=8'b01001101;
   assign rom_data[13524]=8'b00110011;
   assign rom_data[13525]=8'b01001100;
   assign rom_data[13526]=8'b00110011;
   assign rom_data[13527]=8'b01001010;
   assign rom_data[13528]=8'b00110011;
   assign rom_data[13529]=8'b01001001;
   assign rom_data[13530]=8'b00110011;
   assign rom_data[13531]=8'b01000111;
   assign rom_data[13532]=8'b00110011;
   assign rom_data[13533]=8'b01000110;
   assign rom_data[13534]=8'b00110011;
   assign rom_data[13535]=8'b01000101;
   assign rom_data[13536]=8'b00110011;
   assign rom_data[13537]=8'b01000100;
   assign rom_data[13538]=8'b00110011;
   assign rom_data[13539]=8'b01000010;
   assign rom_data[13540]=8'b00110011;
   assign rom_data[13541]=8'b01000001;
   assign rom_data[13542]=8'b00110011;
   assign rom_data[13543]=8'b01000000;
   assign rom_data[13544]=8'b00110011;
   assign rom_data[13545]=8'b00111110;
   assign rom_data[13546]=8'b00110011;
   assign rom_data[13547]=8'b00111101;
   assign rom_data[13548]=8'b00110011;
   assign rom_data[13549]=8'b00111100;
   assign rom_data[13550]=8'b00110011;
   assign rom_data[13551]=8'b00111011;
   assign rom_data[13552]=8'b00110011;
   assign rom_data[13553]=8'b00111010;
   assign rom_data[13554]=8'b00110011;
   assign rom_data[13555]=8'b00111001;
   assign rom_data[13556]=8'b00110011;
   assign rom_data[13557]=8'b00110111;
   assign rom_data[13558]=8'b00110011;
   assign rom_data[13559]=8'b00110110;
   assign rom_data[13560]=8'b00110011;
   assign rom_data[13561]=8'b00110101;
   assign rom_data[13562]=8'b00110010;
   assign rom_data[13563]=8'b00110100;
   assign rom_data[13564]=8'b00110010;
   assign rom_data[13565]=8'b00110011;
   assign rom_data[13566]=8'b00110010;
   assign rom_data[13567]=8'b00110011;
   assign rom_data[13568]=8'b00110010;
   assign rom_data[13569]=8'b00110010;
   assign rom_data[13570]=8'b00110010;
   assign rom_data[13571]=8'b00110001;
   assign rom_data[13572]=8'b00110010;
   assign rom_data[13573]=8'b00110000;
   assign rom_data[13574]=8'b00110010;
   assign rom_data[13575]=8'b00101111;
   assign rom_data[13576]=8'b00110010;
   assign rom_data[13577]=8'b00101111;
   assign rom_data[13578]=8'b00110010;
   assign rom_data[13579]=8'b00101110;
   assign rom_data[13580]=8'b00110010;
   assign rom_data[13581]=8'b00101110;
   assign rom_data[13582]=8'b00110010;
   assign rom_data[13583]=8'b00101101;
   assign rom_data[13584]=8'b00110010;
   assign rom_data[13585]=8'b00101101;
   assign rom_data[13586]=8'b00110010;
   assign rom_data[13587]=8'b00101100;
   assign rom_data[13588]=8'b00110010;
   assign rom_data[13589]=8'b00101100;
   assign rom_data[13590]=8'b00110010;
   assign rom_data[13591]=8'b00101100;
   assign rom_data[13592]=8'b00110010;
   assign rom_data[13593]=8'b00101100;
   assign rom_data[13594]=8'b00110010;
   assign rom_data[13595]=8'b00101100;
   assign rom_data[13596]=8'b00110010;
   assign rom_data[13597]=8'b00101100;
   assign rom_data[13598]=8'b00110010;
   assign rom_data[13599]=8'b00101100;
   assign rom_data[13600]=8'b00110010;
   assign rom_data[13601]=8'b00101101;
   assign rom_data[13602]=8'b00110010;
   assign rom_data[13603]=8'b00101101;
   assign rom_data[13604]=8'b00110010;
   assign rom_data[13605]=8'b00101101;
   assign rom_data[13606]=8'b00110010;
   assign rom_data[13607]=8'b00101110;
   assign rom_data[13608]=8'b00110010;
   assign rom_data[13609]=8'b00101111;
   assign rom_data[13610]=8'b00110010;
   assign rom_data[13611]=8'b00101111;
   assign rom_data[13612]=8'b00110010;
   assign rom_data[13613]=8'b00110000;
   assign rom_data[13614]=8'b00110010;
   assign rom_data[13615]=8'b00110001;
   assign rom_data[13616]=8'b00110010;
   assign rom_data[13617]=8'b00110010;
   assign rom_data[13618]=8'b00110010;
   assign rom_data[13619]=8'b00110010;
   assign rom_data[13620]=8'b00110010;
   assign rom_data[13621]=8'b00110011;
   assign rom_data[13622]=8'b00110010;
   assign rom_data[13623]=8'b00110100;
   assign rom_data[13624]=8'b00110010;
   assign rom_data[13625]=8'b00110101;
   assign rom_data[13626]=8'b00110001;
   assign rom_data[13627]=8'b00110110;
   assign rom_data[13628]=8'b00110001;
   assign rom_data[13629]=8'b00110111;
   assign rom_data[13630]=8'b00110001;
   assign rom_data[13631]=8'b00111001;
   assign rom_data[13632]=8'b00110001;
   assign rom_data[13633]=8'b00111010;
   assign rom_data[13634]=8'b00110001;
   assign rom_data[13635]=8'b00111011;
   assign rom_data[13636]=8'b00110001;
   assign rom_data[13637]=8'b00111100;
   assign rom_data[13638]=8'b00110001;
   assign rom_data[13639]=8'b00111101;
   assign rom_data[13640]=8'b00110001;
   assign rom_data[13641]=8'b00111110;
   assign rom_data[13642]=8'b00110001;
   assign rom_data[13643]=8'b01000000;
   assign rom_data[13644]=8'b00110001;
   assign rom_data[13645]=8'b01000001;
   assign rom_data[13646]=8'b00110001;
   assign rom_data[13647]=8'b01000010;
   assign rom_data[13648]=8'b00110001;
   assign rom_data[13649]=8'b01000100;
   assign rom_data[13650]=8'b00110001;
   assign rom_data[13651]=8'b01000101;
   assign rom_data[13652]=8'b00110001;
   assign rom_data[13653]=8'b01000110;
   assign rom_data[13654]=8'b00110001;
   assign rom_data[13655]=8'b01001000;
   assign rom_data[13656]=8'b00110001;
   assign rom_data[13657]=8'b01001001;
   assign rom_data[13658]=8'b00110001;
   assign rom_data[13659]=8'b01001010;
   assign rom_data[13660]=8'b00110001;
   assign rom_data[13661]=8'b01001100;
   assign rom_data[13662]=8'b00110001;
   assign rom_data[13663]=8'b01001101;
   assign rom_data[13664]=8'b00110001;
   assign rom_data[13665]=8'b01001110;
   assign rom_data[13666]=8'b00110001;
   assign rom_data[13667]=8'b01010000;
   assign rom_data[13668]=8'b00110001;
   assign rom_data[13669]=8'b01010001;
   assign rom_data[13670]=8'b00110001;
   assign rom_data[13671]=8'b01010011;
   assign rom_data[13672]=8'b00110001;
   assign rom_data[13673]=8'b01010100;
   assign rom_data[13674]=8'b00110001;
   assign rom_data[13675]=8'b01010101;
   assign rom_data[13676]=8'b00110001;
   assign rom_data[13677]=8'b01010111;
   assign rom_data[13678]=8'b00110001;
   assign rom_data[13679]=8'b01011000;
   assign rom_data[13680]=8'b00110001;
   assign rom_data[13681]=8'b01011010;
   assign rom_data[13682]=8'b00110001;
   assign rom_data[13683]=8'b01011011;
   assign rom_data[13684]=8'b00110001;
   assign rom_data[13685]=8'b01011100;
   assign rom_data[13686]=8'b00110001;
   assign rom_data[13687]=8'b01011110;
   assign rom_data[13688]=8'b00110001;
   assign rom_data[13689]=8'b01011111;
   assign rom_data[13690]=8'b00110001;
   assign rom_data[13691]=8'b01100001;
   assign rom_data[13692]=8'b00110001;
   assign rom_data[13693]=8'b01100010;
   assign rom_data[13694]=8'b00110001;
   assign rom_data[13695]=8'b01100011;
   assign rom_data[13696]=8'b00110001;
   assign rom_data[13697]=8'b01100101;
   assign rom_data[13698]=8'b00110001;
   assign rom_data[13699]=8'b01100110;
   assign rom_data[13700]=8'b00110001;
   assign rom_data[13701]=8'b01101000;
   assign rom_data[13702]=8'b00110001;
   assign rom_data[13703]=8'b01101001;
   assign rom_data[13704]=8'b00110001;
   assign rom_data[13705]=8'b01101010;
   assign rom_data[13706]=8'b00110001;
   assign rom_data[13707]=8'b01101100;
   assign rom_data[13708]=8'b00110001;
   assign rom_data[13709]=8'b01101101;
   assign rom_data[13710]=8'b00110000;
   assign rom_data[13711]=8'b01101110;
   assign rom_data[13712]=8'b00110000;
   assign rom_data[13713]=8'b01110000;
   assign rom_data[13714]=8'b00110000;
   assign rom_data[13715]=8'b01110001;
   assign rom_data[13716]=8'b00110000;
   assign rom_data[13717]=8'b01110010;
   assign rom_data[13718]=8'b00110000;
   assign rom_data[13719]=8'b01110100;
   assign rom_data[13720]=8'b00110000;
   assign rom_data[13721]=8'b01110101;
   assign rom_data[13722]=8'b00110000;
   assign rom_data[13723]=8'b01110110;
   assign rom_data[13724]=8'b00110000;
   assign rom_data[13725]=8'b01110111;
   assign rom_data[13726]=8'b00110000;
   assign rom_data[13727]=8'b01111001;
   assign rom_data[13728]=8'b00110000;
   assign rom_data[13729]=8'b01111010;
   assign rom_data[13730]=8'b00110000;
   assign rom_data[13731]=8'b01111011;
   assign rom_data[13732]=8'b00110000;
   assign rom_data[13733]=8'b01111100;
   assign rom_data[13734]=8'b00110000;
   assign rom_data[13735]=8'b01111101;
   assign rom_data[13736]=8'b00110000;
   assign rom_data[13737]=8'b01111110;
   assign rom_data[13738]=8'b00110000;
   assign rom_data[13739]=8'b01111111;
   assign rom_data[13740]=8'b00110000;
   assign rom_data[13741]=8'b10000000;
   assign rom_data[13742]=8'b00110000;
   assign rom_data[13743]=8'b10000001;
   assign rom_data[13744]=8'b00110000;
   assign rom_data[13745]=8'b10000010;
   assign rom_data[13746]=8'b00110000;
   assign rom_data[13747]=8'b10000011;
   assign rom_data[13748]=8'b00110000;
   assign rom_data[13749]=8'b10000100;
   assign rom_data[13750]=8'b00110000;
   assign rom_data[13751]=8'b10000101;
   assign rom_data[13752]=8'b00110000;
   assign rom_data[13753]=8'b10000110;
   assign rom_data[13754]=8'b00110000;
   assign rom_data[13755]=8'b10000110;
   assign rom_data[13756]=8'b00110000;
   assign rom_data[13757]=8'b10000111;
   assign rom_data[13758]=8'b00110000;
   assign rom_data[13759]=8'b10001000;
   assign rom_data[13760]=8'b00110000;
   assign rom_data[13761]=8'b10001000;
   assign rom_data[13762]=8'b00110000;
   assign rom_data[13763]=8'b10001001;
   assign rom_data[13764]=8'b00110000;
   assign rom_data[13765]=8'b10001001;
   assign rom_data[13766]=8'b00110000;
   assign rom_data[13767]=8'b10001001;
   assign rom_data[13768]=8'b00110000;
   assign rom_data[13769]=8'b10001010;
   assign rom_data[13770]=8'b00110000;
   assign rom_data[13771]=8'b10001010;
   assign rom_data[13772]=8'b00110000;
   assign rom_data[13773]=8'b10001010;
   assign rom_data[13774]=8'b00110000;
   assign rom_data[13775]=8'b10001010;
   assign rom_data[13776]=8'b00110000;
   assign rom_data[13777]=8'b10001010;
   assign rom_data[13778]=8'b00110000;
   assign rom_data[13779]=8'b10001001;
   assign rom_data[13780]=8'b00101111;
   assign rom_data[13781]=8'b10001001;
   assign rom_data[13782]=8'b00101111;
   assign rom_data[13783]=8'b10001001;
   assign rom_data[13784]=8'b00101111;
   assign rom_data[13785]=8'b10001000;
   assign rom_data[13786]=8'b00101111;
   assign rom_data[13787]=8'b10001000;
   assign rom_data[13788]=8'b00101111;
   assign rom_data[13789]=8'b10000111;
   assign rom_data[13790]=8'b00101111;
   assign rom_data[13791]=8'b10000111;
   assign rom_data[13792]=8'b00101111;
   assign rom_data[13793]=8'b10000110;
   assign rom_data[13794]=8'b00101111;
   assign rom_data[13795]=8'b10000101;
   assign rom_data[13796]=8'b00101111;
   assign rom_data[13797]=8'b10000100;
   assign rom_data[13798]=8'b00101111;
   assign rom_data[13799]=8'b10000011;
   assign rom_data[13800]=8'b00101111;
   assign rom_data[13801]=8'b10000011;
   assign rom_data[13802]=8'b00101111;
   assign rom_data[13803]=8'b10000010;
   assign rom_data[13804]=8'b00101111;
   assign rom_data[13805]=8'b10000001;
   assign rom_data[13806]=8'b00101111;
   assign rom_data[13807]=8'b01111111;
   assign rom_data[13808]=8'b00101111;
   assign rom_data[13809]=8'b01111110;
   assign rom_data[13810]=8'b00101111;
   assign rom_data[13811]=8'b01111101;
   assign rom_data[13812]=8'b00101111;
   assign rom_data[13813]=8'b01111100;
   assign rom_data[13814]=8'b00101111;
   assign rom_data[13815]=8'b01111011;
   assign rom_data[13816]=8'b00101111;
   assign rom_data[13817]=8'b01111010;
   assign rom_data[13818]=8'b00101111;
   assign rom_data[13819]=8'b01111001;
   assign rom_data[13820]=8'b00101111;
   assign rom_data[13821]=8'b01110111;
   assign rom_data[13822]=8'b00101111;
   assign rom_data[13823]=8'b01110110;
   assign rom_data[13824]=8'b00101111;
   assign rom_data[13825]=8'b01110101;
   assign rom_data[13826]=8'b00101111;
   assign rom_data[13827]=8'b01110100;
   assign rom_data[13828]=8'b00101111;
   assign rom_data[13829]=8'b01110010;
   assign rom_data[13830]=8'b00101111;
   assign rom_data[13831]=8'b01110001;
   assign rom_data[13832]=8'b00101111;
   assign rom_data[13833]=8'b01110000;
   assign rom_data[13834]=8'b00101111;
   assign rom_data[13835]=8'b01101110;
   assign rom_data[13836]=8'b00101111;
   assign rom_data[13837]=8'b01101101;
   assign rom_data[13838]=8'b00101111;
   assign rom_data[13839]=8'b01101100;
   assign rom_data[13840]=8'b00101111;
   assign rom_data[13841]=8'b01101010;
   assign rom_data[13842]=8'b00101111;
   assign rom_data[13843]=8'b01101001;
   assign rom_data[13844]=8'b00101111;
   assign rom_data[13845]=8'b01100111;
   assign rom_data[13846]=8'b00101111;
   assign rom_data[13847]=8'b01100110;
   assign rom_data[13848]=8'b00101111;
   assign rom_data[13849]=8'b01100101;
   assign rom_data[13850]=8'b00101111;
   assign rom_data[13851]=8'b01100011;
   assign rom_data[13852]=8'b00101111;
   assign rom_data[13853]=8'b01100010;
   assign rom_data[13854]=8'b00101111;
   assign rom_data[13855]=8'b01100000;
   assign rom_data[13856]=8'b00101110;
   assign rom_data[13857]=8'b01011111;
   assign rom_data[13858]=8'b00101110;
   assign rom_data[13859]=8'b01011110;
   assign rom_data[13860]=8'b00101110;
   assign rom_data[13861]=8'b01011100;
   assign rom_data[13862]=8'b00101110;
   assign rom_data[13863]=8'b01011011;
   assign rom_data[13864]=8'b00101110;
   assign rom_data[13865]=8'b01011001;
   assign rom_data[13866]=8'b00101110;
   assign rom_data[13867]=8'b01011000;
   assign rom_data[13868]=8'b00101110;
   assign rom_data[13869]=8'b01010111;
   assign rom_data[13870]=8'b00101110;
   assign rom_data[13871]=8'b01010101;
   assign rom_data[13872]=8'b00101110;
   assign rom_data[13873]=8'b01010100;
   assign rom_data[13874]=8'b00101110;
   assign rom_data[13875]=8'b01010010;
   assign rom_data[13876]=8'b00101110;
   assign rom_data[13877]=8'b01010001;
   assign rom_data[13878]=8'b00101110;
   assign rom_data[13879]=8'b01010000;
   assign rom_data[13880]=8'b00101110;
   assign rom_data[13881]=8'b01001110;
   assign rom_data[13882]=8'b00101110;
   assign rom_data[13883]=8'b01001101;
   assign rom_data[13884]=8'b00101110;
   assign rom_data[13885]=8'b01001100;
   assign rom_data[13886]=8'b00101110;
   assign rom_data[13887]=8'b01001010;
   assign rom_data[13888]=8'b00101110;
   assign rom_data[13889]=8'b01001001;
   assign rom_data[13890]=8'b00101110;
   assign rom_data[13891]=8'b01000111;
   assign rom_data[13892]=8'b00101110;
   assign rom_data[13893]=8'b01000110;
   assign rom_data[13894]=8'b00101110;
   assign rom_data[13895]=8'b01000101;
   assign rom_data[13896]=8'b00101110;
   assign rom_data[13897]=8'b01000100;
   assign rom_data[13898]=8'b00101110;
   assign rom_data[13899]=8'b01000010;
   assign rom_data[13900]=8'b00101110;
   assign rom_data[13901]=8'b01000001;
   assign rom_data[13902]=8'b00101110;
   assign rom_data[13903]=8'b01000000;
   assign rom_data[13904]=8'b00101110;
   assign rom_data[13905]=8'b00111110;
   assign rom_data[13906]=8'b00101110;
   assign rom_data[13907]=8'b00111101;
   assign rom_data[13908]=8'b00101110;
   assign rom_data[13909]=8'b00111100;
   assign rom_data[13910]=8'b00101110;
   assign rom_data[13911]=8'b00111011;
   assign rom_data[13912]=8'b00101110;
   assign rom_data[13913]=8'b00111010;
   assign rom_data[13914]=8'b00101110;
   assign rom_data[13915]=8'b00111001;
   assign rom_data[13916]=8'b00101110;
   assign rom_data[13917]=8'b00110111;
   assign rom_data[13918]=8'b00101110;
   assign rom_data[13919]=8'b00110110;
   assign rom_data[13920]=8'b00101110;
   assign rom_data[13921]=8'b00110101;
   assign rom_data[13922]=8'b00101110;
   assign rom_data[13923]=8'b00110100;
   assign rom_data[13924]=8'b00101110;
   assign rom_data[13925]=8'b00110011;
   assign rom_data[13926]=8'b00101110;
   assign rom_data[13927]=8'b00110011;
   assign rom_data[13928]=8'b00101110;
   assign rom_data[13929]=8'b00110010;
   assign rom_data[13930]=8'b00101110;
   assign rom_data[13931]=8'b00110001;
   assign rom_data[13932]=8'b00101110;
   assign rom_data[13933]=8'b00110000;
   assign rom_data[13934]=8'b00101101;
   assign rom_data[13935]=8'b00101111;
   assign rom_data[13936]=8'b00101101;
   assign rom_data[13937]=8'b00101111;
   assign rom_data[13938]=8'b00101101;
   assign rom_data[13939]=8'b00101110;
   assign rom_data[13940]=8'b00101101;
   assign rom_data[13941]=8'b00101110;
   assign rom_data[13942]=8'b00101101;
   assign rom_data[13943]=8'b00101101;
   assign rom_data[13944]=8'b00101101;
   assign rom_data[13945]=8'b00101101;
   assign rom_data[13946]=8'b00101101;
   assign rom_data[13947]=8'b00101100;
   assign rom_data[13948]=8'b00101101;
   assign rom_data[13949]=8'b00101100;
   assign rom_data[13950]=8'b00101101;
   assign rom_data[13951]=8'b00101100;
   assign rom_data[13952]=8'b00101101;
   assign rom_data[13953]=8'b00101100;
   assign rom_data[13954]=8'b00101101;
   assign rom_data[13955]=8'b00101100;
   assign rom_data[13956]=8'b00101101;
   assign rom_data[13957]=8'b00101100;
   assign rom_data[13958]=8'b00101101;
   assign rom_data[13959]=8'b00101100;
   assign rom_data[13960]=8'b00101101;
   assign rom_data[13961]=8'b00101101;
   assign rom_data[13962]=8'b00101101;
   assign rom_data[13963]=8'b00101101;
   assign rom_data[13964]=8'b00101101;
   assign rom_data[13965]=8'b00101101;
   assign rom_data[13966]=8'b00101101;
   assign rom_data[13967]=8'b00101110;
   assign rom_data[13968]=8'b00101101;
   assign rom_data[13969]=8'b00101111;
   assign rom_data[13970]=8'b00101101;
   assign rom_data[13971]=8'b00101111;
   assign rom_data[13972]=8'b00101101;
   assign rom_data[13973]=8'b00110000;
   assign rom_data[13974]=8'b00101101;
   assign rom_data[13975]=8'b00110001;
   assign rom_data[13976]=8'b00101101;
   assign rom_data[13977]=8'b00110010;
   assign rom_data[13978]=8'b00101101;
   assign rom_data[13979]=8'b00110010;
   assign rom_data[13980]=8'b00101101;
   assign rom_data[13981]=8'b00110011;
   assign rom_data[13982]=8'b00101101;
   assign rom_data[13983]=8'b00110100;
   assign rom_data[13984]=8'b00101101;
   assign rom_data[13985]=8'b00110101;
   assign rom_data[13986]=8'b00101101;
   assign rom_data[13987]=8'b00110110;
   assign rom_data[13988]=8'b00101101;
   assign rom_data[13989]=8'b00110111;
   assign rom_data[13990]=8'b00101101;
   assign rom_data[13991]=8'b00111001;
   assign rom_data[13992]=8'b00101101;
   assign rom_data[13993]=8'b00111010;
   assign rom_data[13994]=8'b00101101;
   assign rom_data[13995]=8'b00111011;
   assign rom_data[13996]=8'b00101101;
   assign rom_data[13997]=8'b00111100;
   assign rom_data[13998]=8'b00101101;
   assign rom_data[13999]=8'b00111101;
   assign rom_data[14000]=8'b00101101;
   assign rom_data[14001]=8'b00111110;
   assign rom_data[14002]=8'b00101101;
   assign rom_data[14003]=8'b01000000;
   assign rom_data[14004]=8'b00101101;
   assign rom_data[14005]=8'b01000001;
   assign rom_data[14006]=8'b00101101;
   assign rom_data[14007]=8'b01000010;
   assign rom_data[14008]=8'b00101101;
   assign rom_data[14009]=8'b01000100;
   assign rom_data[14010]=8'b00101100;
   assign rom_data[14011]=8'b01000101;
   assign rom_data[14012]=8'b00101100;
   assign rom_data[14013]=8'b01000110;
   assign rom_data[14014]=8'b00101100;
   assign rom_data[14015]=8'b01001000;
   assign rom_data[14016]=8'b00101100;
   assign rom_data[14017]=8'b01001001;
   assign rom_data[14018]=8'b00101100;
   assign rom_data[14019]=8'b01001010;
   assign rom_data[14020]=8'b00101100;
   assign rom_data[14021]=8'b01001100;
   assign rom_data[14022]=8'b00101100;
   assign rom_data[14023]=8'b01001101;
   assign rom_data[14024]=8'b00101100;
   assign rom_data[14025]=8'b01001110;
   assign rom_data[14026]=8'b00101100;
   assign rom_data[14027]=8'b01010000;
   assign rom_data[14028]=8'b00101100;
   assign rom_data[14029]=8'b01010001;
   assign rom_data[14030]=8'b00101100;
   assign rom_data[14031]=8'b01010011;
   assign rom_data[14032]=8'b00101100;
   assign rom_data[14033]=8'b01010100;
   assign rom_data[14034]=8'b00101100;
   assign rom_data[14035]=8'b01010101;
   assign rom_data[14036]=8'b00101100;
   assign rom_data[14037]=8'b01010111;
   assign rom_data[14038]=8'b00101100;
   assign rom_data[14039]=8'b01011000;
   assign rom_data[14040]=8'b00101100;
   assign rom_data[14041]=8'b01011010;

   // assign rom_data[17716]=8'b01001011;
   // assign rom_data[17717]=8'b10000111;
   // assign rom_data[17718]=8'b01001011;
   // assign rom_data[17719]=8'b10001000;
   // assign rom_data[17720]=8'b01001011;
   // assign rom_data[17721]=8'b10001000;
   // assign rom_data[17722]=8'b01001011;
   // assign rom_data[17723]=8'b10001001;
   // assign rom_data[17724]=8'b01001011;
   // assign rom_data[17725]=8'b10001001;
   // assign rom_data[17726]=8'b01001011;
   // assign rom_data[17727]=8'b10001001;
   // assign rom_data[17728]=8'b01001011;
   // assign rom_data[17729]=8'b10001010;
   // assign rom_data[17730]=8'b01001011;
   // assign rom_data[17731]=8'b10001010;
   // assign rom_data[17732]=8'b01001011;
   // assign rom_data[17733]=8'b10001010;
   // assign rom_data[17734]=8'b01001011;
   // assign rom_data[17735]=8'b10001010;
   // assign rom_data[17736]=8'b01001011;
   // assign rom_data[17737]=8'b10001010;
   // assign rom_data[17738]=8'b01001011;
   // assign rom_data[17739]=8'b10001001;
   // assign rom_data[17740]=8'b01001011;
   // assign rom_data[17741]=8'b10001001;
   // assign rom_data[17742]=8'b01001011;
   // assign rom_data[17743]=8'b10001001;
   // assign rom_data[17744]=8'b01001011;
   // assign rom_data[17745]=8'b10001000;
   // assign rom_data[17746]=8'b01001011;
   // assign rom_data[17747]=8'b10001000;
   // assign rom_data[17748]=8'b01001011;
   // assign rom_data[17749]=8'b10000111;
   // assign rom_data[17750]=8'b01001011;
   // assign rom_data[17751]=8'b10000111;
   // assign rom_data[17752]=8'b01001011;
   // assign rom_data[17753]=8'b10000110;
   // assign rom_data[17754]=8'b01001011;
   // assign rom_data[17755]=8'b10000101;
   // assign rom_data[17756]=8'b01001011;
   // assign rom_data[17757]=8'b10000100;
   // assign rom_data[17758]=8'b01001011;
   // assign rom_data[17759]=8'b10000011;
   // assign rom_data[17760]=8'b01001011;
   // assign rom_data[17761]=8'b10000010;
   // assign rom_data[17762]=8'b01001011;
   // assign rom_data[17763]=8'b10000010;
   // assign rom_data[17764]=8'b01001011;
   // assign rom_data[17765]=8'b10000001;
   // assign rom_data[17766]=8'b01001011;
   // assign rom_data[17767]=8'b01111111;
   // assign rom_data[17768]=8'b01001011;
   // assign rom_data[17769]=8'b01111110;
   // assign rom_data[17770]=8'b01001011;
   // assign rom_data[17771]=8'b01111101;
   // assign rom_data[17772]=8'b01001011;
   // assign rom_data[17773]=8'b01111100;
   // assign rom_data[17774]=8'b01001011;
   // assign rom_data[17775]=8'b01111011;
   // assign rom_data[17776]=8'b01001011;
   // assign rom_data[17777]=8'b01111010;
   // assign rom_data[17778]=8'b01001011;
   // assign rom_data[17779]=8'b01111001;
   // assign rom_data[17780]=8'b01001011;
   // assign rom_data[17781]=8'b01110111;
   // assign rom_data[17782]=8'b01001011;
   // assign rom_data[17783]=8'b01110110;
   // assign rom_data[17784]=8'b01001011;
   // assign rom_data[17785]=8'b01110101;
   // assign rom_data[17786]=8'b01001010;
   // assign rom_data[17787]=8'b01110100;
   // assign rom_data[17788]=8'b01001010;
   // assign rom_data[17789]=8'b01110010;
   // assign rom_data[17790]=8'b01001010;
   // assign rom_data[17791]=8'b01110001;
   // assign rom_data[17792]=8'b01001010;
   // assign rom_data[17793]=8'b01110000;
   // assign rom_data[17794]=8'b01001010;
   // assign rom_data[17795]=8'b01101110;
   // assign rom_data[17796]=8'b01001010;
   // assign rom_data[17797]=8'b01101101;
   // assign rom_data[17798]=8'b01001010;
   // assign rom_data[17799]=8'b01101100;
   // assign rom_data[17800]=8'b01001010;
   // assign rom_data[17801]=8'b01101010;
   // assign rom_data[17802]=8'b01001010;
   // assign rom_data[17803]=8'b01101001;
   // assign rom_data[17804]=8'b01001010;
   // assign rom_data[17805]=8'b01100111;
   // assign rom_data[17806]=8'b01001010;
   // assign rom_data[17807]=8'b01100110;
   // assign rom_data[17808]=8'b01001010;
   // assign rom_data[17809]=8'b01100101;
   // assign rom_data[17810]=8'b01001010;
   // assign rom_data[17811]=8'b01100011;
   // assign rom_data[17812]=8'b01001010;
   // assign rom_data[17813]=8'b01100010;
   // assign rom_data[17814]=8'b01001010;
   // assign rom_data[17815]=8'b01100000;
   // assign rom_data[17816]=8'b01001010;
   // assign rom_data[17817]=8'b01011111;
   // assign rom_data[17818]=8'b01001010;
   // assign rom_data[17819]=8'b01011110;
   // assign rom_data[17820]=8'b01001010;
   // assign rom_data[17821]=8'b01011100;
   // assign rom_data[17822]=8'b01001010;
   // assign rom_data[17823]=8'b01011011;
   // assign rom_data[17824]=8'b01001010;
   // assign rom_data[17825]=8'b01011001;
   // assign rom_data[17826]=8'b01001010;
   // assign rom_data[17827]=8'b01011000;
   // assign rom_data[17828]=8'b01001010;
   // assign rom_data[17829]=8'b01010111;
   // assign rom_data[17830]=8'b01001010;
   // assign rom_data[17831]=8'b01010101;
   // assign rom_data[17832]=8'b01001010;
   // assign rom_data[17833]=8'b01010100;
   // assign rom_data[17834]=8'b01001010;
   // assign rom_data[17835]=8'b01010010;
   // assign rom_data[17836]=8'b01001010;
   // assign rom_data[17837]=8'b01010001;
   // assign rom_data[17838]=8'b01001010;
   // assign rom_data[17839]=8'b01010000;
   // assign rom_data[17840]=8'b01001010;
   // assign rom_data[17841]=8'b01001110;
   // assign rom_data[17842]=8'b01001010;
   // assign rom_data[17843]=8'b01001101;
   // assign rom_data[17844]=8'b01001010;
   // assign rom_data[17845]=8'b01001100;
   // assign rom_data[17846]=8'b01001010;
   // assign rom_data[17847]=8'b01001010;
   // assign rom_data[17848]=8'b01001010;
   // assign rom_data[17849]=8'b01001001;
   // assign rom_data[17850]=8'b01001010;
   // assign rom_data[17851]=8'b01000111;
   // assign rom_data[17852]=8'b01001010;
   // assign rom_data[17853]=8'b01000110;
   // assign rom_data[17854]=8'b01001010;
   // assign rom_data[17855]=8'b01000101;
   // assign rom_data[17856]=8'b01001010;
   // assign rom_data[17857]=8'b01000100;
   // assign rom_data[17858]=8'b01001010;
   // assign rom_data[17859]=8'b01000010;
   // assign rom_data[17860]=8'b01001010;
   // assign rom_data[17861]=8'b01000001;
   // assign rom_data[17862]=8'b01001010;
   // assign rom_data[17863]=8'b01000000;
   // assign rom_data[17864]=8'b01001010;
   // assign rom_data[17865]=8'b00111110;
   // assign rom_data[17866]=8'b01001010;
   // assign rom_data[17867]=8'b00111101;
   // assign rom_data[17868]=8'b01001010;
   // assign rom_data[17869]=8'b00111100;
   // assign rom_data[17870]=8'b01001010;
   // assign rom_data[17871]=8'b00111011;
   // assign rom_data[17872]=8'b01001010;
   // assign rom_data[17873]=8'b00111010;
   // assign rom_data[17874]=8'b01001010;
   // assign rom_data[17875]=8'b00111001;
   // assign rom_data[17876]=8'b01001010;
   // assign rom_data[17877]=8'b00110111;
   // assign rom_data[17878]=8'b01001010;
   // assign rom_data[17879]=8'b00110110;
   // assign rom_data[17880]=8'b01001010;
   // assign rom_data[17881]=8'b00110101;
   // assign rom_data[17882]=8'b01001010;
   // assign rom_data[17883]=8'b00110100;
   // assign rom_data[17884]=8'b01001010;
   // assign rom_data[17885]=8'b00110011;
   // assign rom_data[17886]=8'b01001010;
   // assign rom_data[17887]=8'b00110010;
   // assign rom_data[17888]=8'b01001010;
   // assign rom_data[17889]=8'b00110010;
   // assign rom_data[17890]=8'b01001010;
   // assign rom_data[17891]=8'b00110001;
   // assign rom_data[17892]=8'b01001010;
   // assign rom_data[17893]=8'b00110000;
   // assign rom_data[17894]=8'b01001010;
   // assign rom_data[17895]=8'b00101111;
   // assign rom_data[17896]=8'b01001010;
   // assign rom_data[17897]=8'b00101111;
   // assign rom_data[17898]=8'b01001010;
   // assign rom_data[17899]=8'b00101110;
   // assign rom_data[17900]=8'b01001010;
   // assign rom_data[17901]=8'b00101110;
   // assign rom_data[17902]=8'b01001010;
   // assign rom_data[17903]=8'b00101101;
   // assign rom_data[17904]=8'b01001001;
   // assign rom_data[17905]=8'b00101101;
   // assign rom_data[17906]=8'b01001001;
   // assign rom_data[17907]=8'b00101100;
   // assign rom_data[17908]=8'b01001001;
   // assign rom_data[17909]=8'b00101100;
   // assign rom_data[17910]=8'b01001001;
   // assign rom_data[17911]=8'b00101100;
   // assign rom_data[17912]=8'b01001001;
   // assign rom_data[17913]=8'b00101100;
   // assign rom_data[17914]=8'b01001001;
   // assign rom_data[17915]=8'b00101100;
   // assign rom_data[17916]=8'b01001001;
   // assign rom_data[17917]=8'b00101100;
   // assign rom_data[17918]=8'b01001001;
   // assign rom_data[17919]=8'b00101100;
   // assign rom_data[17920]=8'b01001001;
   // assign rom_data[17921]=8'b00101101;
   // assign rom_data[17922]=8'b01001001;
   // assign rom_data[17923]=8'b00101101;
   // assign rom_data[17924]=8'b01001001;
   // assign rom_data[17925]=8'b00101101;
   // assign rom_data[17926]=8'b01001001;
   // assign rom_data[17927]=8'b00101110;
   // assign rom_data[17928]=8'b01001001;
   // assign rom_data[17929]=8'b00101111;
   // assign rom_data[17930]=8'b01001001;
   // assign rom_data[17931]=8'b00101111;
   // assign rom_data[17932]=8'b01001001;
   // assign rom_data[17933]=8'b00110000;
   // assign rom_data[17934]=8'b01001001;
   // assign rom_data[17935]=8'b00110001;
   // assign rom_data[17936]=8'b01001001;
   // assign rom_data[17937]=8'b00110010;
   // assign rom_data[17938]=8'b01001001;
   // assign rom_data[17939]=8'b00110010;
   // assign rom_data[17940]=8'b01001001;
   // assign rom_data[17941]=8'b00110011;
   // assign rom_data[17942]=8'b01001001;
   // assign rom_data[17943]=8'b00110100;
   // assign rom_data[17944]=8'b01001001;
   // assign rom_data[17945]=8'b00110101;
   // assign rom_data[17946]=8'b01001001;
   // assign rom_data[17947]=8'b00110110;
   // assign rom_data[17948]=8'b01001001;
   // assign rom_data[17949]=8'b00110111;
   // assign rom_data[17950]=8'b01001001;
   // assign rom_data[17951]=8'b00111001;
   // assign rom_data[17952]=8'b01001001;
   // assign rom_data[17953]=8'b00111010;
   // assign rom_data[17954]=8'b01001001;
   // assign rom_data[17955]=8'b00111011;
   // assign rom_data[17956]=8'b01001001;
   // assign rom_data[17957]=8'b00111100;
   // assign rom_data[17958]=8'b01001001;
   // assign rom_data[17959]=8'b00111101;
   // assign rom_data[17960]=8'b01001001;
   // assign rom_data[17961]=8'b00111110;
   // assign rom_data[17962]=8'b01001001;
   // assign rom_data[17963]=8'b01000000;
   // assign rom_data[17964]=8'b01001001;
   // assign rom_data[17965]=8'b01000001;
   // assign rom_data[17966]=8'b01001001;
   // assign rom_data[17967]=8'b01000010;
   // assign rom_data[17968]=8'b01001001;
   // assign rom_data[17969]=8'b01000100;
   // assign rom_data[17970]=8'b01001001;
   // assign rom_data[17971]=8'b01000101;
   // assign rom_data[17972]=8'b01001001;
   // assign rom_data[17973]=8'b01000110;
   // assign rom_data[17974]=8'b01001001;
   // assign rom_data[17975]=8'b01001000;
   // assign rom_data[17976]=8'b01001001;
   // assign rom_data[17977]=8'b01001001;
   // assign rom_data[17978]=8'b01001001;
   // assign rom_data[17979]=8'b01001010;
   // assign rom_data[17980]=8'b01001001;
   // assign rom_data[17981]=8'b01001100;
   // assign rom_data[17982]=8'b01001001;
   // assign rom_data[17983]=8'b01001101;
   // assign rom_data[17984]=8'b01001001;
   // assign rom_data[17985]=8'b01001110;
   // assign rom_data[17986]=8'b01001001;
   // assign rom_data[17987]=8'b01010000;
   // assign rom_data[17988]=8'b01001001;
   // assign rom_data[17989]=8'b01010001;
   // assign rom_data[17990]=8'b01001001;
   // assign rom_data[17991]=8'b01010011;
   // assign rom_data[17992]=8'b01001001;
   // assign rom_data[17993]=8'b01010100;
   // assign rom_data[17994]=8'b01001001;
   // assign rom_data[17995]=8'b01010101;
   // assign rom_data[17996]=8'b01001001;
   // assign rom_data[17997]=8'b01010111;
   // assign rom_data[17998]=8'b01001001;
   // assign rom_data[17999]=8'b01011000;
   // assign rom_data[18000]=8'b01001001;
   // assign rom_data[18001]=8'b01011010;
   // assign rom_data[18002]=8'b01001001;
   // assign rom_data[18003]=8'b01011011;
   // assign rom_data[18004]=8'b01001001;
   // assign rom_data[18005]=8'b01011100;
   // assign rom_data[18006]=8'b01001001;
   // assign rom_data[18007]=8'b01011110;
   // assign rom_data[18008]=8'b01001001;
   // assign rom_data[18009]=8'b01011111;
   // assign rom_data[18010]=8'b01001001;
   // assign rom_data[18011]=8'b01100001;
   // assign rom_data[18012]=8'b01001001;
   // assign rom_data[18013]=8'b01100010;
   // assign rom_data[18014]=8'b01001001;
   // assign rom_data[18015]=8'b01100011;
   // assign rom_data[18016]=8'b01001001;
   // assign rom_data[18017]=8'b01100101;
   // assign rom_data[18018]=8'b01001001;
   // assign rom_data[18019]=8'b01100110;
   // assign rom_data[18020]=8'b01001000;
   // assign rom_data[18021]=8'b01101000;
   // assign rom_data[18022]=8'b01001000;
   // assign rom_data[18023]=8'b01101001;
   // assign rom_data[18024]=8'b01001000;
   // assign rom_data[18025]=8'b01101010;
   // assign rom_data[18026]=8'b01001000;
   // assign rom_data[18027]=8'b01101100;
   // assign rom_data[18028]=8'b01001000;
   // assign rom_data[18029]=8'b01101101;
   // assign rom_data[18030]=8'b01001000;
   // assign rom_data[18031]=8'b01101110;
   // assign rom_data[18032]=8'b01001000;
   // assign rom_data[18033]=8'b01110000;
   // assign rom_data[18034]=8'b01001000;
   // assign rom_data[18035]=8'b01110001;
   // assign rom_data[18036]=8'b01001000;
   // assign rom_data[18037]=8'b01110010;
   // assign rom_data[18038]=8'b01001000;
   // assign rom_data[18039]=8'b01110100;
   // assign rom_data[18040]=8'b01001000;
   // assign rom_data[18041]=8'b01110101;
   // assign rom_data[18042]=8'b01001000;
   // assign rom_data[18043]=8'b01110110;
   // assign rom_data[18044]=8'b01001000;
   // assign rom_data[18045]=8'b01110111;
   // assign rom_data[18046]=8'b01001000;
   // assign rom_data[18047]=8'b01111001;
   // assign rom_data[18048]=8'b01001000;
   // assign rom_data[18049]=8'b01111010;
   // assign rom_data[18050]=8'b01001000;
   // assign rom_data[18051]=8'b01111011;
   // assign rom_data[18052]=8'b01001000;
   // assign rom_data[18053]=8'b01111100;
   // assign rom_data[18054]=8'b01001000;
   // assign rom_data[18055]=8'b01111101;
   // assign rom_data[18056]=8'b01001000;
   // assign rom_data[18057]=8'b01111110;
   // assign rom_data[18058]=8'b01001000;
   // assign rom_data[18059]=8'b01111111;
   // assign rom_data[18060]=8'b01001000;
   // assign rom_data[18061]=8'b10000000;
   // assign rom_data[18062]=8'b01001000;
   // assign rom_data[18063]=8'b10000001;
   // assign rom_data[18064]=8'b01001000;
   // assign rom_data[18065]=8'b10000010;
   // assign rom_data[18066]=8'b01001000;
   // assign rom_data[18067]=8'b10000011;
   // assign rom_data[18068]=8'b01001000;
   // assign rom_data[18069]=8'b10000100;
   // assign rom_data[18070]=8'b01001000;
   // assign rom_data[18071]=8'b10000101;
   // assign rom_data[18072]=8'b01001000;
   // assign rom_data[18073]=8'b10000110;
   // assign rom_data[18074]=8'b01001000;
   // assign rom_data[18075]=8'b10000110;
   // assign rom_data[18076]=8'b01001000;
   // assign rom_data[18077]=8'b10000111;
   // assign rom_data[18078]=8'b01001000;
   // assign rom_data[18079]=8'b10001000;
   // assign rom_data[18080]=8'b01001000;
   // assign rom_data[18081]=8'b10001000;
   // assign rom_data[18082]=8'b01001000;
   // assign rom_data[18083]=8'b10001001;
   // assign rom_data[18084]=8'b01001000;
   // assign rom_data[18085]=8'b10001001;
   // assign rom_data[18086]=8'b01001000;
   // assign rom_data[18087]=8'b10001001;
   // assign rom_data[18088]=8'b01001000;
   // assign rom_data[18089]=8'b10001010;
   // assign rom_data[18090]=8'b01001000;
   // assign rom_data[18091]=8'b10001010;
   // assign rom_data[18092]=8'b01001000;
   // assign rom_data[18093]=8'b10001010;
   // assign rom_data[18094]=8'b01001000;
   // assign rom_data[18095]=8'b10001010;
   // assign rom_data[18096]=8'b01001000;
   // assign rom_data[18097]=8'b10001010;
   // assign rom_data[18098]=8'b01001000;
   // assign rom_data[18099]=8'b10001001;
   // assign rom_data[18100]=8'b01001000;
   // assign rom_data[18101]=8'b10001001;
   // assign rom_data[18102]=8'b01001000;
   // assign rom_data[18103]=8'b10001001;
   // assign rom_data[18104]=8'b01001000;
   // assign rom_data[18105]=8'b10001000;
   // assign rom_data[18106]=8'b01001000;
   // assign rom_data[18107]=8'b10001000;
   // assign rom_data[18108]=8'b01001000;
   // assign rom_data[18109]=8'b10000111;
   // assign rom_data[18110]=8'b01001000;
   // assign rom_data[18111]=8'b10000111;
   // assign rom_data[18112]=8'b01001000;
   // assign rom_data[18113]=8'b10000110;
   // assign rom_data[18114]=8'b01001000;
   // assign rom_data[18115]=8'b10000101;
   // assign rom_data[18116]=8'b01001000;
   // assign rom_data[18117]=8'b10000100;
   // assign rom_data[18118]=8'b01001000;
   // assign rom_data[18119]=8'b10000011;
   // assign rom_data[18120]=8'b01001000;
   // assign rom_data[18121]=8'b10000010;
   // assign rom_data[18122]=8'b01001000;
   // assign rom_data[18123]=8'b10000010;
   // assign rom_data[18124]=8'b01001000;
   // assign rom_data[18125]=8'b10000001;
   // assign rom_data[18126]=8'b01000111;
   // assign rom_data[18127]=8'b01111111;
   // assign rom_data[18128]=8'b01000111;
   // assign rom_data[18129]=8'b01111110;
   // assign rom_data[18130]=8'b01000111;
   // assign rom_data[18131]=8'b01111101;
   // assign rom_data[18132]=8'b01000111;
   // assign rom_data[18133]=8'b01111100;
   // assign rom_data[18134]=8'b01000111;
   // assign rom_data[18135]=8'b01111011;
   // assign rom_data[18136]=8'b01000111;
   // assign rom_data[18137]=8'b01111010;
   // assign rom_data[18138]=8'b01000111;
   // assign rom_data[18139]=8'b01111001;
   // assign rom_data[18140]=8'b01000111;
   // assign rom_data[18141]=8'b01110111;
   // assign rom_data[18142]=8'b01000111;
   // assign rom_data[18143]=8'b01110110;
   // assign rom_data[18144]=8'b01000111;
   // assign rom_data[18145]=8'b01110101;
   // assign rom_data[18146]=8'b01000111;
   // assign rom_data[18147]=8'b01110100;
   // assign rom_data[18148]=8'b01000111;
   // assign rom_data[18149]=8'b01110010;
   // assign rom_data[18150]=8'b01000111;
   // assign rom_data[18151]=8'b01110001;
   // assign rom_data[18152]=8'b01000111;
   // assign rom_data[18153]=8'b01110000;
   // assign rom_data[18154]=8'b01000111;
   // assign rom_data[18155]=8'b01101110;
   // assign rom_data[18156]=8'b01000111;
   // assign rom_data[18157]=8'b01101101;
   // assign rom_data[18158]=8'b01000111;
   // assign rom_data[18159]=8'b01101100;
   // assign rom_data[18160]=8'b01000111;
   // assign rom_data[18161]=8'b01101010;
   // assign rom_data[18162]=8'b01000111;
   // assign rom_data[18163]=8'b01101001;
   // assign rom_data[18164]=8'b01000111;
   // assign rom_data[18165]=8'b01100111;
   // assign rom_data[18166]=8'b01000111;
   // assign rom_data[18167]=8'b01100110;
   // assign rom_data[18168]=8'b01000111;
   // assign rom_data[18169]=8'b01100101;
   // assign rom_data[18170]=8'b01000111;
   // assign rom_data[18171]=8'b01100011;
   // assign rom_data[18172]=8'b01000111;
   // assign rom_data[18173]=8'b01100010;
   // assign rom_data[18174]=8'b01000111;
   // assign rom_data[18175]=8'b01100000;
   // assign rom_data[18176]=8'b01000111;
   // assign rom_data[18177]=8'b01011111;
   // assign rom_data[18178]=8'b01000111;
   // assign rom_data[18179]=8'b01011110;
   // assign rom_data[18180]=8'b01000111;
   // assign rom_data[18181]=8'b01011100;
   // assign rom_data[18182]=8'b01000111;
   // assign rom_data[18183]=8'b01011011;
   // assign rom_data[18184]=8'b01000111;
   // assign rom_data[18185]=8'b01011001;
   // assign rom_data[18186]=8'b01000111;
   // assign rom_data[18187]=8'b01011000;
   // assign rom_data[18188]=8'b01000111;
   // assign rom_data[18189]=8'b01010111;
   // assign rom_data[18190]=8'b01000111;
   // assign rom_data[18191]=8'b01010101;
   // assign rom_data[18192]=8'b01000111;
   // assign rom_data[18193]=8'b01010100;
   // assign rom_data[18194]=8'b01000111;
   // assign rom_data[18195]=8'b01010010;
   // assign rom_data[18196]=8'b01000111;
   // assign rom_data[18197]=8'b01010001;
   // assign rom_data[18198]=8'b01000111;
   // assign rom_data[18199]=8'b01010000;
   // assign rom_data[18200]=8'b01000111;
   // assign rom_data[18201]=8'b01001110;
   // assign rom_data[18202]=8'b01000111;
   // assign rom_data[18203]=8'b01001101;
   // assign rom_data[18204]=8'b01000111;
   // assign rom_data[18205]=8'b01001100;
   // assign rom_data[18206]=8'b01000111;
   // assign rom_data[18207]=8'b01001010;
   // assign rom_data[18208]=8'b01000111;
   // assign rom_data[18209]=8'b01001001;
   // assign rom_data[18210]=8'b01000111;
   // assign rom_data[18211]=8'b01000111;
   // assign rom_data[18212]=8'b01000111;
   // assign rom_data[18213]=8'b01000110;
   // assign rom_data[18214]=8'b01000111;
   // assign rom_data[18215]=8'b01000101;
   // assign rom_data[18216]=8'b01000111;
   // assign rom_data[18217]=8'b01000100;
   // assign rom_data[18218]=8'b01000111;
   // assign rom_data[18219]=8'b01000010;
   // assign rom_data[18220]=8'b01000111;
   // assign rom_data[18221]=8'b01000001;
   // assign rom_data[18222]=8'b01000111;
   // assign rom_data[18223]=8'b01000000;
   // assign rom_data[18224]=8'b01000111;
   // assign rom_data[18225]=8'b00111110;
   // assign rom_data[18226]=8'b01000111;
   // assign rom_data[18227]=8'b00111101;
   // assign rom_data[18228]=8'b01000111;
   // assign rom_data[18229]=8'b00111100;
   // assign rom_data[18230]=8'b01000111;
   // assign rom_data[18231]=8'b00111011;
   // assign rom_data[18232]=8'b01000111;
   // assign rom_data[18233]=8'b00111010;
   // assign rom_data[18234]=8'b01000111;
   // assign rom_data[18235]=8'b00111001;
   // assign rom_data[18236]=8'b01000111;
   // assign rom_data[18237]=8'b00110111;
   // assign rom_data[18238]=8'b01000111;
   // assign rom_data[18239]=8'b00110110;
   // assign rom_data[18240]=8'b01000111;
   // assign rom_data[18241]=8'b00110101;
   // assign rom_data[18242]=8'b01000111;
   // assign rom_data[18243]=8'b00110100;
   // assign rom_data[18244]=8'b01000111;
   // assign rom_data[18245]=8'b00110011;
   // assign rom_data[18246]=8'b01000111;
   // assign rom_data[18247]=8'b00110010;
   // assign rom_data[18248]=8'b01000110;
   // assign rom_data[18249]=8'b00110010;
   // assign rom_data[18250]=8'b01000110;
   // assign rom_data[18251]=8'b00110001;
   // assign rom_data[18252]=8'b01000110;
   // assign rom_data[18253]=8'b00110000;
   // assign rom_data[18254]=8'b01000110;
   // assign rom_data[18255]=8'b00101111;
   // assign rom_data[18256]=8'b01000110;
   // assign rom_data[18257]=8'b00101111;
   // assign rom_data[18258]=8'b01000110;
   // assign rom_data[18259]=8'b00101110;
   // assign rom_data[18260]=8'b01000110;
   // assign rom_data[18261]=8'b00101110;
   // assign rom_data[18262]=8'b01000110;
   // assign rom_data[18263]=8'b00101101;
   // assign rom_data[18264]=8'b01000110;
   // assign rom_data[18265]=8'b00101101;
   // assign rom_data[18266]=8'b01000110;
   // assign rom_data[18267]=8'b00101100;
   // assign rom_data[18268]=8'b01000110;
   // assign rom_data[18269]=8'b00101100;
   // assign rom_data[18270]=8'b01000110;
   // assign rom_data[18271]=8'b00101100;
   // assign rom_data[18272]=8'b01000110;
   // assign rom_data[18273]=8'b00101100;
   // assign rom_data[18274]=8'b01000110;
   // assign rom_data[18275]=8'b00101100;
   // assign rom_data[18276]=8'b01000110;
   // assign rom_data[18277]=8'b00101100;
   // assign rom_data[18278]=8'b01000110;
   // assign rom_data[18279]=8'b00101100;
   // assign rom_data[18280]=8'b01000110;
   // assign rom_data[18281]=8'b00101101;
   // assign rom_data[18282]=8'b01000110;
   // assign rom_data[18283]=8'b00101101;
   // assign rom_data[18284]=8'b01000110;
   // assign rom_data[18285]=8'b00101101;
   // assign rom_data[18286]=8'b01000110;
   // assign rom_data[18287]=8'b00101110;
   // assign rom_data[18288]=8'b01000110;
   // assign rom_data[18289]=8'b00101111;
   // assign rom_data[18290]=8'b01000110;
   // assign rom_data[18291]=8'b00101111;
   // assign rom_data[18292]=8'b01000110;
   // assign rom_data[18293]=8'b00110000;
   // assign rom_data[18294]=8'b01000110;
   // assign rom_data[18295]=8'b00110001;
   // assign rom_data[18296]=8'b01000110;
   // assign rom_data[18297]=8'b00110010;
   // assign rom_data[18298]=8'b01000110;
   // assign rom_data[18299]=8'b00110010;
   // assign rom_data[18300]=8'b01000110;
   // assign rom_data[18301]=8'b00110011;
   // assign rom_data[18302]=8'b01000110;
   // assign rom_data[18303]=8'b00110100;
   // assign rom_data[18304]=8'b01000110;
   // assign rom_data[18305]=8'b00110101;
   // assign rom_data[18306]=8'b01000110;
   // assign rom_data[18307]=8'b00110110;
   // assign rom_data[18308]=8'b01000110;
   // assign rom_data[18309]=8'b00110111;
   // assign rom_data[18310]=8'b01000110;
   // assign rom_data[18311]=8'b00111001;
   // assign rom_data[18312]=8'b01000110;
   // assign rom_data[18313]=8'b00111010;
   // assign rom_data[18314]=8'b01000110;
   // assign rom_data[18315]=8'b00111011;
   // assign rom_data[18316]=8'b01000110;
   // assign rom_data[18317]=8'b00111100;
   // assign rom_data[18318]=8'b01000110;
   // assign rom_data[18319]=8'b00111101;
   // assign rom_data[18320]=8'b01000110;
   // assign rom_data[18321]=8'b00111110;
   // assign rom_data[18322]=8'b01000110;
   // assign rom_data[18323]=8'b01000000;
   // assign rom_data[18324]=8'b01000110;
   // assign rom_data[18325]=8'b01000001;
   // assign rom_data[18326]=8'b01000110;
   // assign rom_data[18327]=8'b01000010;
   // assign rom_data[18328]=8'b01000110;
   // assign rom_data[18329]=8'b01000100;
   // assign rom_data[18330]=8'b01000110;
   // assign rom_data[18331]=8'b01000101;
   // assign rom_data[18332]=8'b01000110;
   // assign rom_data[18333]=8'b01000110;
   // assign rom_data[18334]=8'b01000110;
   // assign rom_data[18335]=8'b01001000;
   // assign rom_data[18336]=8'b01000110;
   // assign rom_data[18337]=8'b01001001;
   // assign rom_data[18338]=8'b01000110;
   // assign rom_data[18339]=8'b01001010;
   // assign rom_data[18340]=8'b01000110;
   // assign rom_data[18341]=8'b01001100;
   // assign rom_data[18342]=8'b01000110;
   // assign rom_data[18343]=8'b01001101;
   // assign rom_data[18344]=8'b01000110;
   // assign rom_data[18345]=8'b01001110;
   // assign rom_data[18346]=8'b01000110;
   // assign rom_data[18347]=8'b01010000;
   // assign rom_data[18348]=8'b01000110;
   // assign rom_data[18349]=8'b01010001;
   // assign rom_data[18350]=8'b01000110;
   // assign rom_data[18351]=8'b01010011;
   // assign rom_data[18352]=8'b01000110;
   // assign rom_data[18353]=8'b01010100;
   // assign rom_data[18354]=8'b01000110;
   // assign rom_data[18355]=8'b01010101;
   // assign rom_data[18356]=8'b01000101;
   // assign rom_data[18357]=8'b01010111;
   // assign rom_data[18358]=8'b01000101;
   // assign rom_data[18359]=8'b01011000;
   // assign rom_data[18360]=8'b01000101;
   // assign rom_data[18361]=8'b01011010;
   // assign rom_data[18362]=8'b01000101;
   // assign rom_data[18363]=8'b01011011;
   // assign rom_data[18364]=8'b01000101;
   // assign rom_data[18365]=8'b01011100;
   // assign rom_data[18366]=8'b01000101;
   // assign rom_data[18367]=8'b01011110;
   // assign rom_data[18368]=8'b01000101;
   // assign rom_data[18369]=8'b01011111;
   // assign rom_data[18370]=8'b01000101;
   // assign rom_data[18371]=8'b01100001;
   // assign rom_data[18372]=8'b01000101;
   // assign rom_data[18373]=8'b01100010;
   // assign rom_data[18374]=8'b01000101;
   // assign rom_data[18375]=8'b01100011;
   // assign rom_data[18376]=8'b01000101;
   // assign rom_data[18377]=8'b01100101;
   // assign rom_data[18378]=8'b01000101;
   // assign rom_data[18379]=8'b01100110;
   // assign rom_data[18380]=8'b01000101;
   // assign rom_data[18381]=8'b01101000;
   // assign rom_data[18382]=8'b01000101;
   // assign rom_data[18383]=8'b01101001;
   // assign rom_data[18384]=8'b01000101;
   // assign rom_data[18385]=8'b01101010;
   // assign rom_data[18386]=8'b01000101;
   // assign rom_data[18387]=8'b01101100;
   // assign rom_data[18388]=8'b01000101;
   // assign rom_data[18389]=8'b01101101;
   // assign rom_data[18390]=8'b01000101;
   // assign rom_data[18391]=8'b01101110;
   // assign rom_data[18392]=8'b01000101;
   // assign rom_data[18393]=8'b01110000;
   // assign rom_data[18394]=8'b01000101;
   // assign rom_data[18395]=8'b01110001;
   // assign rom_data[18396]=8'b01000101;
   // assign rom_data[18397]=8'b01110010;
   // assign rom_data[18398]=8'b01000101;
   // assign rom_data[18399]=8'b01110100;
   // assign rom_data[18400]=8'b01000101;
   // assign rom_data[18401]=8'b01110101;
   // assign rom_data[18402]=8'b01000101;
   // assign rom_data[18403]=8'b01110110;
   // assign rom_data[18404]=8'b01000101;
   // assign rom_data[18405]=8'b01110111;
   // assign rom_data[18406]=8'b01000101;
   // assign rom_data[18407]=8'b01111001;
   // assign rom_data[18408]=8'b01000101;
   // assign rom_data[18409]=8'b01111010;
   // assign rom_data[18410]=8'b01000101;
   // assign rom_data[18411]=8'b01111011;
   // assign rom_data[18412]=8'b01000101;
   // assign rom_data[18413]=8'b01111100;
   // assign rom_data[18414]=8'b01000101;
   // assign rom_data[18415]=8'b01111101;
   // assign rom_data[18416]=8'b01000101;
   // assign rom_data[18417]=8'b01111110;
   // assign rom_data[18418]=8'b01000101;
   // assign rom_data[18419]=8'b01111111;
   // assign rom_data[18420]=8'b01000101;
   // assign rom_data[18421]=8'b10000000;
   // assign rom_data[18422]=8'b01000101;
   // assign rom_data[18423]=8'b10000001;
   // assign rom_data[18424]=8'b01000101;
   // assign rom_data[18425]=8'b10000010;
   // assign rom_data[18426]=8'b01000101;
   // assign rom_data[18427]=8'b10000011;
   // assign rom_data[18428]=8'b01000101;
   // assign rom_data[18429]=8'b10000100;
   // assign rom_data[18430]=8'b01000101;
   // assign rom_data[18431]=8'b10000101;
   // assign rom_data[18432]=8'b01000101;
   // assign rom_data[18433]=8'b10000110;
   // assign rom_data[18434]=8'b01000101;
   // assign rom_data[18435]=8'b10000110;
   // assign rom_data[18436]=8'b01000101;
   // assign rom_data[18437]=8'b10000111;
   // assign rom_data[18438]=8'b01000101;
   // assign rom_data[18439]=8'b10001000;
   // assign rom_data[18440]=8'b01000101;
   // assign rom_data[18441]=8'b10001000;
   // assign rom_data[18442]=8'b01000101;
   // assign rom_data[18443]=8'b10001001;
   // assign rom_data[18444]=8'b01000101;
   // assign rom_data[18445]=8'b10001001;
   // assign rom_data[18446]=8'b01000101;
   // assign rom_data[18447]=8'b10001001;
   // assign rom_data[18448]=8'b01000101;
   // assign rom_data[18449]=8'b10001010;
   // assign rom_data[18450]=8'b01000101;
   // assign rom_data[18451]=8'b10001010;
   // assign rom_data[18452]=8'b01000101;
   // assign rom_data[18453]=8'b10001010;
   // assign rom_data[18454]=8'b01000101;
   // assign rom_data[18455]=8'b10001010;
   // assign rom_data[18456]=8'b01000101;
   // assign rom_data[18457]=8'b10001010;
   // assign rom_data[18458]=8'b01000101;
   // assign rom_data[18459]=8'b10001001;
   // assign rom_data[18460]=8'b01000101;
   // assign rom_data[18461]=8'b10001001;
   // assign rom_data[18462]=8'b01000101;
   // assign rom_data[18463]=8'b10001001;
   // assign rom_data[18464]=8'b01000101;
   // assign rom_data[18465]=8'b10001000;
   // assign rom_data[18466]=8'b01000100;
   // assign rom_data[18467]=8'b10001000;
   // assign rom_data[18468]=8'b01000100;
   // assign rom_data[18469]=8'b10000111;
   // assign rom_data[18470]=8'b01000100;
   // assign rom_data[18471]=8'b10000111;
   // assign rom_data[18472]=8'b01000100;
   // assign rom_data[18473]=8'b10000110;
   // assign rom_data[18474]=8'b01000100;
   // assign rom_data[18475]=8'b10000101;
   // assign rom_data[18476]=8'b01000100;
   // assign rom_data[18477]=8'b10000100;
   // assign rom_data[18478]=8'b01000100;
   // assign rom_data[18479]=8'b10000011;
   // assign rom_data[18480]=8'b01000100;
   // assign rom_data[18481]=8'b10000010;
   // assign rom_data[18482]=8'b01000100;
   // assign rom_data[18483]=8'b10000010;
   // assign rom_data[18484]=8'b01000100;
   // assign rom_data[18485]=8'b10000001;
   // assign rom_data[18486]=8'b01000100;
   // assign rom_data[18487]=8'b01111111;
   // assign rom_data[18488]=8'b01000100;
   // assign rom_data[18489]=8'b01111110;
   // assign rom_data[18490]=8'b01000100;
   // assign rom_data[18491]=8'b01111101;
   // assign rom_data[18492]=8'b01000100;
   // assign rom_data[18493]=8'b01111100;
   // assign rom_data[18494]=8'b01000100;
   // assign rom_data[18495]=8'b01111011;
   // assign rom_data[18496]=8'b01000100;
   // assign rom_data[18497]=8'b01111010;
   // assign rom_data[18498]=8'b01000100;
   // assign rom_data[18499]=8'b01111001;
   // assign rom_data[18500]=8'b01000100;
   // assign rom_data[18501]=8'b01110111;
   // assign rom_data[18502]=8'b01000100;
   // assign rom_data[18503]=8'b01110110;
   // assign rom_data[18504]=8'b01000100;
   // assign rom_data[18505]=8'b01110101;
   // assign rom_data[18506]=8'b01000100;
   // assign rom_data[18507]=8'b01110100;
   // assign rom_data[18508]=8'b01000100;
   // assign rom_data[18509]=8'b01110010;
   // assign rom_data[18510]=8'b01000100;
   // assign rom_data[18511]=8'b01110001;
   // assign rom_data[18512]=8'b01000100;
   // assign rom_data[18513]=8'b01110000;
   // assign rom_data[18514]=8'b01000100;
   // assign rom_data[18515]=8'b01101110;
   // assign rom_data[18516]=8'b01000100;
   // assign rom_data[18517]=8'b01101101;
   // assign rom_data[18518]=8'b01000100;
   // assign rom_data[18519]=8'b01101100;
   // assign rom_data[18520]=8'b01000100;
   // assign rom_data[18521]=8'b01101010;
   // assign rom_data[18522]=8'b01000100;
   // assign rom_data[18523]=8'b01101001;
   // assign rom_data[18524]=8'b01000100;
   // assign rom_data[18525]=8'b01100111;
   // assign rom_data[18526]=8'b01000100;
   // assign rom_data[18527]=8'b01100110;
   // assign rom_data[18528]=8'b01000100;
   // assign rom_data[18529]=8'b01100101;
   // assign rom_data[18530]=8'b01000100;
   // assign rom_data[18531]=8'b01100011;
   // assign rom_data[18532]=8'b01000100;
   // assign rom_data[18533]=8'b01100010;
   // assign rom_data[18534]=8'b01000100;
   // assign rom_data[18535]=8'b01100000;
   // assign rom_data[18536]=8'b01000100;
   // assign rom_data[18537]=8'b01011111;
   // assign rom_data[18538]=8'b01000100;
   // assign rom_data[18539]=8'b01011110;
   // assign rom_data[18540]=8'b01000100;
   // assign rom_data[18541]=8'b01011100;
   // assign rom_data[18542]=8'b01000100;
   // assign rom_data[18543]=8'b01011011;
   // assign rom_data[18544]=8'b01000100;
   // assign rom_data[18545]=8'b01011001;
   // assign rom_data[18546]=8'b01000100;
   // assign rom_data[18547]=8'b01011000;
   // assign rom_data[18548]=8'b01000100;
   // assign rom_data[18549]=8'b01010111;
   // assign rom_data[18550]=8'b01000100;
   // assign rom_data[18551]=8'b01010101;
   // assign rom_data[18552]=8'b01000100;
   // assign rom_data[18553]=8'b01010100;
   // assign rom_data[18554]=8'b01000100;
   // assign rom_data[18555]=8'b01010010;
   // assign rom_data[18556]=8'b01000100;
   // assign rom_data[18557]=8'b01010001;
   // assign rom_data[18558]=8'b01000100;
   // assign rom_data[18559]=8'b01010000;
   // assign rom_data[18560]=8'b01000100;
   // assign rom_data[18561]=8'b01001110;
   // assign rom_data[18562]=8'b01000100;
   // assign rom_data[18563]=8'b01001101;
   // assign rom_data[18564]=8'b01000100;
   // assign rom_data[18565]=8'b01001100;
   // assign rom_data[18566]=8'b01000100;
   // assign rom_data[18567]=8'b01001010;
   // assign rom_data[18568]=8'b01000100;
   // assign rom_data[18569]=8'b01001001;
   // assign rom_data[18570]=8'b01000100;
   // assign rom_data[18571]=8'b01000111;
   // assign rom_data[18572]=8'b01000100;
   // assign rom_data[18573]=8'b01000110;
   // assign rom_data[18574]=8'b01000100;
   // assign rom_data[18575]=8'b01000101;
   // assign rom_data[18576]=8'b01000100;
   // assign rom_data[18577]=8'b01000100;
   // assign rom_data[18578]=8'b01000100;
   // assign rom_data[18579]=8'b01000010;
   // assign rom_data[18580]=8'b01000100;
   // assign rom_data[18581]=8'b01000001;
   // assign rom_data[18582]=8'b01000100;
   // assign rom_data[18583]=8'b01000000;
   // assign rom_data[18584]=8'b01000100;
   // assign rom_data[18585]=8'b00111110;
   // assign rom_data[18586]=8'b01000100;
   // assign rom_data[18587]=8'b00111101;
   // assign rom_data[18588]=8'b01000011;
   // assign rom_data[18589]=8'b00111100;
   // assign rom_data[18590]=8'b01000011;
   // assign rom_data[18591]=8'b00111011;
   // assign rom_data[18592]=8'b01000011;
   // assign rom_data[18593]=8'b00111010;
   // assign rom_data[18594]=8'b01000011;
   // assign rom_data[18595]=8'b00111001;
   // assign rom_data[18596]=8'b01000011;
   // assign rom_data[18597]=8'b00110111;
   // assign rom_data[18598]=8'b01000011;
   // assign rom_data[18599]=8'b00110110;
   // assign rom_data[18600]=8'b01000011;
   // assign rom_data[18601]=8'b00110101;
   // assign rom_data[18602]=8'b01000011;
   // assign rom_data[18603]=8'b00110100;
   // assign rom_data[18604]=8'b01000011;
   // assign rom_data[18605]=8'b00110011;
   // assign rom_data[18606]=8'b01000011;
   // assign rom_data[18607]=8'b00110010;
   // assign rom_data[18608]=8'b01000011;
   // assign rom_data[18609]=8'b00110010;
   // assign rom_data[18610]=8'b01000011;
   // assign rom_data[18611]=8'b00110001;
   // assign rom_data[18612]=8'b01000011;
   // assign rom_data[18613]=8'b00110000;
   // assign rom_data[18614]=8'b01000011;
   // assign rom_data[18615]=8'b00101111;
   // assign rom_data[18616]=8'b01000011;
   // assign rom_data[18617]=8'b00101111;
   // assign rom_data[18618]=8'b01000011;
   // assign rom_data[18619]=8'b00101110;
   // assign rom_data[18620]=8'b01000011;
   // assign rom_data[18621]=8'b00101110;
   // assign rom_data[18622]=8'b01000011;
   // assign rom_data[18623]=8'b00101101;
   // assign rom_data[18624]=8'b01000011;
   // assign rom_data[18625]=8'b00101101;
   // assign rom_data[18626]=8'b01000011;
   // assign rom_data[18627]=8'b00101100;
   // assign rom_data[18628]=8'b01000011;
   // assign rom_data[18629]=8'b00101100;
   // assign rom_data[18630]=8'b01000011;
   // assign rom_data[18631]=8'b00101100;
   // assign rom_data[18632]=8'b01000011;
   // assign rom_data[18633]=8'b00101100;
   // assign rom_data[18634]=8'b01000011;
   // assign rom_data[18635]=8'b00101100;
   // assign rom_data[18636]=8'b01000011;
   // assign rom_data[18637]=8'b00101100;
   // assign rom_data[18638]=8'b01000011;
   // assign rom_data[18639]=8'b00101100;
   // assign rom_data[18640]=8'b01000011;
   // assign rom_data[18641]=8'b00101101;
   // assign rom_data[18642]=8'b01000011;
   // assign rom_data[18643]=8'b00101101;
   // assign rom_data[18644]=8'b01000011;
   // assign rom_data[18645]=8'b00101101;
   // assign rom_data[18646]=8'b01000011;
   // assign rom_data[18647]=8'b00101110;
   // assign rom_data[18648]=8'b01000011;
   // assign rom_data[18649]=8'b00101111;
   // assign rom_data[18650]=8'b01000011;
   // assign rom_data[18651]=8'b00101111;
   // assign rom_data[18652]=8'b01000011;
   // assign rom_data[18653]=8'b00110000;
   // assign rom_data[18654]=8'b01000011;
   // assign rom_data[18655]=8'b00110001;
   // assign rom_data[18656]=8'b01000011;
   // assign rom_data[18657]=8'b00110010;
   // assign rom_data[18658]=8'b01000011;
   // assign rom_data[18659]=8'b00110010;
   // assign rom_data[18660]=8'b01000011;
   // assign rom_data[18661]=8'b00110011;
   // assign rom_data[18662]=8'b01000011;
   // assign rom_data[18663]=8'b00110100;
   // assign rom_data[18664]=8'b01000011;
   // assign rom_data[18665]=8'b00110101;
   // assign rom_data[18666]=8'b01000011;
   // assign rom_data[18667]=8'b00110110;
   // assign rom_data[18668]=8'b01000011;
   // assign rom_data[18669]=8'b00110111;
   // assign rom_data[18670]=8'b01000011;
   // assign rom_data[18671]=8'b00111001;
   // assign rom_data[18672]=8'b01000011;
   // assign rom_data[18673]=8'b00111010;
   // assign rom_data[18674]=8'b01000011;
   // assign rom_data[18675]=8'b00111011;
   // assign rom_data[18676]=8'b01000011;
   // assign rom_data[18677]=8'b00111100;
   // assign rom_data[18678]=8'b01000011;
   // assign rom_data[18679]=8'b00111101;
   // assign rom_data[18680]=8'b01000011;
   // assign rom_data[18681]=8'b00111110;
   // assign rom_data[18682]=8'b01000011;
   // assign rom_data[18683]=8'b01000000;
   // assign rom_data[18684]=8'b01000011;
   // assign rom_data[18685]=8'b01000001;
   // assign rom_data[18686]=8'b01000011;
   // assign rom_data[18687]=8'b01000010;
   // assign rom_data[18688]=8'b01000011;
   // assign rom_data[18689]=8'b01000100;
   // assign rom_data[18690]=8'b01000011;
   // assign rom_data[18691]=8'b01000101;
   // assign rom_data[18692]=8'b01000010;
   // assign rom_data[18693]=8'b01000110;
   // assign rom_data[18694]=8'b01000010;
   // assign rom_data[18695]=8'b01001000;
   // assign rom_data[18696]=8'b01000010;
   // assign rom_data[18697]=8'b01001001;
   // assign rom_data[18698]=8'b01000010;
   // assign rom_data[18699]=8'b01001010;
   // assign rom_data[18700]=8'b01000010;
   // assign rom_data[18701]=8'b01001100;
   // assign rom_data[18702]=8'b01000010;
   // assign rom_data[18703]=8'b01001101;
   // assign rom_data[18704]=8'b01000010;
   // assign rom_data[18705]=8'b01001110;
   // assign rom_data[18706]=8'b01000010;
   // assign rom_data[18707]=8'b01010000;
   // assign rom_data[18708]=8'b01000010;
   // assign rom_data[18709]=8'b01010001;
   // assign rom_data[18710]=8'b01000010;
   // assign rom_data[18711]=8'b01010011;
   // assign rom_data[18712]=8'b01000010;
   // assign rom_data[18713]=8'b01010100;
   // assign rom_data[18714]=8'b01000010;
   // assign rom_data[18715]=8'b01010101;
   // assign rom_data[18716]=8'b01000010;
   // assign rom_data[18717]=8'b01010111;
   // assign rom_data[18718]=8'b01000010;
   // assign rom_data[18719]=8'b01011000;
   // assign rom_data[18720]=8'b01000010;
   // assign rom_data[18721]=8'b01011010;
   // assign rom_data[18722]=8'b01000010;
   // assign rom_data[18723]=8'b01011011;
   // assign rom_data[18724]=8'b01000010;
   // assign rom_data[18725]=8'b01011100;
   // assign rom_data[18726]=8'b01000010;
   // assign rom_data[18727]=8'b01011110;
   // assign rom_data[18728]=8'b01000010;
   // assign rom_data[18729]=8'b01011111;
   // assign rom_data[18730]=8'b01000010;
   // assign rom_data[18731]=8'b01100001;
   // assign rom_data[18732]=8'b01000010;
   // assign rom_data[18733]=8'b01100010;
   // assign rom_data[18734]=8'b01000010;
   // assign rom_data[18735]=8'b01100011;
   // assign rom_data[18736]=8'b01000010;
   // assign rom_data[18737]=8'b01100101;
   // assign rom_data[18738]=8'b01000010;
   // assign rom_data[18739]=8'b01100110;
   // assign rom_data[18740]=8'b01000010;
   // assign rom_data[18741]=8'b01101000;
   // assign rom_data[18742]=8'b01000010;
   // assign rom_data[18743]=8'b01101001;
   // assign rom_data[18744]=8'b01000010;
   // assign rom_data[18745]=8'b01101010;
   // assign rom_data[18746]=8'b01000010;
   // assign rom_data[18747]=8'b01101100;
   // assign rom_data[18748]=8'b01000010;
   // assign rom_data[18749]=8'b01101101;
   // assign rom_data[18750]=8'b01000010;
   // assign rom_data[18751]=8'b01101110;
   // assign rom_data[18752]=8'b01000010;
   // assign rom_data[18753]=8'b01110000;
   // assign rom_data[18754]=8'b01000010;
   // assign rom_data[18755]=8'b01110001;
   // assign rom_data[18756]=8'b01000010;
   // assign rom_data[18757]=8'b01110010;
   // assign rom_data[18758]=8'b01000010;
   // assign rom_data[18759]=8'b01110100;
   // assign rom_data[18760]=8'b01000010;
   // assign rom_data[18761]=8'b01110101;
   // assign rom_data[18762]=8'b01000010;
   // assign rom_data[18763]=8'b01110110;
   // assign rom_data[18764]=8'b01000010;
   // assign rom_data[18765]=8'b01110111;
   // assign rom_data[18766]=8'b01000010;
   // assign rom_data[18767]=8'b01111001;
   // assign rom_data[18768]=8'b01000010;
   // assign rom_data[18769]=8'b01111010;
   // assign rom_data[18770]=8'b01000010;
   // assign rom_data[18771]=8'b01111011;
   // assign rom_data[18772]=8'b01000010;
   // assign rom_data[18773]=8'b01111100;
   // assign rom_data[18774]=8'b01000010;
   // assign rom_data[18775]=8'b01111101;
   // assign rom_data[18776]=8'b01000010;
   // assign rom_data[18777]=8'b01111110;
   // assign rom_data[18778]=8'b01000010;
   // assign rom_data[18779]=8'b01111111;
   // assign rom_data[18780]=8'b01000010;
   // assign rom_data[18781]=8'b10000000;
   // assign rom_data[18782]=8'b01000010;
   // assign rom_data[18783]=8'b10000001;
   // assign rom_data[18784]=8'b01000010;
   // assign rom_data[18785]=8'b10000010;
   // assign rom_data[18786]=8'b01000010;
   // assign rom_data[18787]=8'b10000011;
   // assign rom_data[18788]=8'b01000010;
   // assign rom_data[18789]=8'b10000100;
   // assign rom_data[18790]=8'b01000010;
   // assign rom_data[18791]=8'b10000101;
   // assign rom_data[18792]=8'b01000010;
   // assign rom_data[18793]=8'b10000110;
   // assign rom_data[18794]=8'b01000010;
   // assign rom_data[18795]=8'b10000110;
   // assign rom_data[18796]=8'b01000010;
   // assign rom_data[18797]=8'b10000111;
   // assign rom_data[18798]=8'b01000010;
   // assign rom_data[18799]=8'b10001000;
   // assign rom_data[18800]=8'b01000010;
   // assign rom_data[18801]=8'b10001000;
   // assign rom_data[18802]=8'b01000010;
   // assign rom_data[18803]=8'b10001001;
   // assign rom_data[18804]=8'b01000010;
   // assign rom_data[18805]=8'b10001001;
   // assign rom_data[18806]=8'b01000010;
   // assign rom_data[18807]=8'b10001001;
   // assign rom_data[18808]=8'b01000010;
   // assign rom_data[18809]=8'b10001010;
   // assign rom_data[18810]=8'b01000001;
   // assign rom_data[18811]=8'b10001010;
   // assign rom_data[18812]=8'b01000001;
   // assign rom_data[18813]=8'b10001010;
   // assign rom_data[18814]=8'b01000001;
   // assign rom_data[18815]=8'b10001010;
   // assign rom_data[18816]=8'b01000001;
   // assign rom_data[18817]=8'b10001010;
   // assign rom_data[18818]=8'b01000001;
   // assign rom_data[18819]=8'b10001001;
   // assign rom_data[18820]=8'b01000001;
   // assign rom_data[18821]=8'b10001001;
   // assign rom_data[18822]=8'b01000001;
   // assign rom_data[18823]=8'b10001001;
   // assign rom_data[18824]=8'b01000001;
   // assign rom_data[18825]=8'b10001000;
   // assign rom_data[18826]=8'b01000001;
   // assign rom_data[18827]=8'b10001000;
   // assign rom_data[18828]=8'b01000001;
   // assign rom_data[18829]=8'b10000111;
   // assign rom_data[18830]=8'b01000001;
   // assign rom_data[18831]=8'b10000111;
   // assign rom_data[18832]=8'b01000001;
   // assign rom_data[18833]=8'b10000110;
   // assign rom_data[18834]=8'b01000001;
   // assign rom_data[18835]=8'b10000101;
   // assign rom_data[18836]=8'b01000001;
   // assign rom_data[18837]=8'b10000100;
   // assign rom_data[18838]=8'b01000001;
   // assign rom_data[18839]=8'b10000011;
   // assign rom_data[18840]=8'b01000001;
   // assign rom_data[18841]=8'b10000010;
   // assign rom_data[18842]=8'b01000001;
   // assign rom_data[18843]=8'b10000010;
   // assign rom_data[18844]=8'b01000001;
   // assign rom_data[18845]=8'b10000001;
   // assign rom_data[18846]=8'b01000001;
   // assign rom_data[18847]=8'b01111111;
   // assign rom_data[18848]=8'b01000001;
   // assign rom_data[18849]=8'b01111110;
   // assign rom_data[18850]=8'b01000001;
   // assign rom_data[18851]=8'b01111101;
   // assign rom_data[18852]=8'b01000001;
   // assign rom_data[18853]=8'b01111100;
   // assign rom_data[18854]=8'b01000001;
   // assign rom_data[18855]=8'b01111011;
   // assign rom_data[18856]=8'b01000001;
   // assign rom_data[18857]=8'b01111010;
   // assign rom_data[18858]=8'b01000001;
   // assign rom_data[18859]=8'b01111001;
   // assign rom_data[18860]=8'b01000001;
   // assign rom_data[18861]=8'b01110111;
   // assign rom_data[18862]=8'b01000001;
   // assign rom_data[18863]=8'b01110110;
   // assign rom_data[18864]=8'b01000001;
   // assign rom_data[18865]=8'b01110101;
   // assign rom_data[18866]=8'b01000001;
   // assign rom_data[18867]=8'b01110100;
   // assign rom_data[18868]=8'b01000001;
   // assign rom_data[18869]=8'b01110010;
   // assign rom_data[18870]=8'b01000001;
   // assign rom_data[18871]=8'b01110001;
   // assign rom_data[18872]=8'b01000001;
   // assign rom_data[18873]=8'b01110000;
   // assign rom_data[18874]=8'b01000001;
   // assign rom_data[18875]=8'b01101110;
   // assign rom_data[18876]=8'b01000001;
   // assign rom_data[18877]=8'b01101101;
   // assign rom_data[18878]=8'b01000001;
   // assign rom_data[18879]=8'b01101100;
   // assign rom_data[18880]=8'b01000001;
   // assign rom_data[18881]=8'b01101010;
   // assign rom_data[18882]=8'b01000001;
   // assign rom_data[18883]=8'b01101001;
   // assign rom_data[18884]=8'b01000001;
   // assign rom_data[18885]=8'b01100111;
   // assign rom_data[18886]=8'b01000001;
   // assign rom_data[18887]=8'b01100110;
   // assign rom_data[18888]=8'b01000001;
   // assign rom_data[18889]=8'b01100101;
   // assign rom_data[18890]=8'b01000001;
   // assign rom_data[18891]=8'b01100011;
   // assign rom_data[18892]=8'b01000001;
   // assign rom_data[18893]=8'b01100010;
   // assign rom_data[18894]=8'b01000001;
   // assign rom_data[18895]=8'b01100000;
   // assign rom_data[18896]=8'b01000001;
   // assign rom_data[18897]=8'b01011111;
   // assign rom_data[18898]=8'b01000001;
   // assign rom_data[18899]=8'b01011110;
   // assign rom_data[18900]=8'b01000001;
   // assign rom_data[18901]=8'b01011100;
   // assign rom_data[18902]=8'b01000001;
   // assign rom_data[18903]=8'b01011011;
   // assign rom_data[18904]=8'b01000001;
   // assign rom_data[18905]=8'b01011001;
   // assign rom_data[18906]=8'b01000001;
   // assign rom_data[18907]=8'b01011000;
   // assign rom_data[18908]=8'b01000001;
   // assign rom_data[18909]=8'b01010111;
   // assign rom_data[18910]=8'b01000001;
   // assign rom_data[18911]=8'b01010101;
   // assign rom_data[18912]=8'b01000001;
   // assign rom_data[18913]=8'b01010100;
   // assign rom_data[18914]=8'b01000001;
   // assign rom_data[18915]=8'b01010010;
   // assign rom_data[18916]=8'b01000001;
   // assign rom_data[18917]=8'b01010001;
   // assign rom_data[18918]=8'b01000001;
   // assign rom_data[18919]=8'b01010000;
   // assign rom_data[18920]=8'b01000001;
   // assign rom_data[18921]=8'b01001110;
   // assign rom_data[18922]=8'b01000001;
   // assign rom_data[18923]=8'b01001101;
   // assign rom_data[18924]=8'b01000001;
   // assign rom_data[18925]=8'b01001100;
   // assign rom_data[18926]=8'b01000000;
   // assign rom_data[18927]=8'b01001010;
   // assign rom_data[18928]=8'b01000000;
   // assign rom_data[18929]=8'b01001001;
   // assign rom_data[18930]=8'b01000000;
   // assign rom_data[18931]=8'b01000111;
   // assign rom_data[18932]=8'b01000000;
   // assign rom_data[18933]=8'b01000110;
   // assign rom_data[18934]=8'b01000000;
   // assign rom_data[18935]=8'b01000101;
   // assign rom_data[18936]=8'b01000000;
   // assign rom_data[18937]=8'b01000100;
   // assign rom_data[18938]=8'b01000000;
   // assign rom_data[18939]=8'b01000010;
   // assign rom_data[18940]=8'b01000000;
   // assign rom_data[18941]=8'b01000001;
   // assign rom_data[18942]=8'b01000000;
   // assign rom_data[18943]=8'b01000000;
   // assign rom_data[18944]=8'b01000000;
   // assign rom_data[18945]=8'b00111110;
   // assign rom_data[18946]=8'b01000000;
   // assign rom_data[18947]=8'b00111101;
   // assign rom_data[18948]=8'b01000000;
   // assign rom_data[18949]=8'b00111100;
   // assign rom_data[18950]=8'b01000000;
   // assign rom_data[18951]=8'b00111011;
   // assign rom_data[18952]=8'b01000000;
   // assign rom_data[18953]=8'b00111010;
   // assign rom_data[18954]=8'b01000000;
   // assign rom_data[18955]=8'b00111001;
   // assign rom_data[18956]=8'b01000000;
   // assign rom_data[18957]=8'b00110111;
   // assign rom_data[18958]=8'b01000000;
   // assign rom_data[18959]=8'b00110110;
   // assign rom_data[18960]=8'b01000000;
   // assign rom_data[18961]=8'b00110101;
   // assign rom_data[18962]=8'b01000000;
   // assign rom_data[18963]=8'b00110100;
   // assign rom_data[18964]=8'b01000000;
   // assign rom_data[18965]=8'b00110011;
   // assign rom_data[18966]=8'b01000000;
   // assign rom_data[18967]=8'b00110010;
   // assign rom_data[18968]=8'b01000000;
   // assign rom_data[18969]=8'b00110010;
   // assign rom_data[18970]=8'b01000000;
   // assign rom_data[18971]=8'b00110001;
   // assign rom_data[18972]=8'b01000000;
   // assign rom_data[18973]=8'b00110000;
   // assign rom_data[18974]=8'b01000000;
   // assign rom_data[18975]=8'b00101111;
   // assign rom_data[18976]=8'b01000000;
   // assign rom_data[18977]=8'b00101111;
   // assign rom_data[18978]=8'b01000000;
   // assign rom_data[18979]=8'b00101110;
   // assign rom_data[18980]=8'b01000000;
   // assign rom_data[18981]=8'b00101110;
   // assign rom_data[18982]=8'b01000000;
   // assign rom_data[18983]=8'b00101101;
   // assign rom_data[18984]=8'b01000000;
   // assign rom_data[18985]=8'b00101101;
   // assign rom_data[18986]=8'b01000000;
   // assign rom_data[18987]=8'b00101100;
   // assign rom_data[18988]=8'b01000000;
   // assign rom_data[18989]=8'b00101100;
   // assign rom_data[18990]=8'b01000000;
   // assign rom_data[18991]=8'b00101100;
   // assign rom_data[18992]=8'b01000000;
   // assign rom_data[18993]=8'b00101100;
   // assign rom_data[18994]=8'b01000000;
   // assign rom_data[18995]=8'b00101100;
   // assign rom_data[18996]=8'b01000000;
   // assign rom_data[18997]=8'b00101100;
   // assign rom_data[18998]=8'b01000000;
   // assign rom_data[18999]=8'b00101100;
   // assign rom_data[19000]=8'b01000000;
   // assign rom_data[19001]=8'b00101101;
   // assign rom_data[19002]=8'b01000000;
   // assign rom_data[19003]=8'b00101101;
   // assign rom_data[19004]=8'b01000000;
   // assign rom_data[19005]=8'b00101101;
   // assign rom_data[19006]=8'b01000000;
   // assign rom_data[19007]=8'b00101110;
   // assign rom_data[19008]=8'b01000000;
   // assign rom_data[19009]=8'b00101111;
   // assign rom_data[19010]=8'b01000000;
   // assign rom_data[19011]=8'b00101111;
   // assign rom_data[19012]=8'b01000000;
   // assign rom_data[19013]=8'b00110000;
   // assign rom_data[19014]=8'b01000000;
   // assign rom_data[19015]=8'b00110001;
   // assign rom_data[19016]=8'b01000000;
   // assign rom_data[19017]=8'b00110010;
   // assign rom_data[19018]=8'b01000000;
   // assign rom_data[19019]=8'b00110010;
   // assign rom_data[19020]=8'b01000000;
   // assign rom_data[19021]=8'b00110011;
   // assign rom_data[19022]=8'b01000000;
   // assign rom_data[19023]=8'b00110100;
   // assign rom_data[19024]=8'b01000000;
   // assign rom_data[19025]=8'b00110101;
   // assign rom_data[19026]=8'b01000000;
   // assign rom_data[19027]=8'b00110110;
   // assign rom_data[19028]=8'b01000000;
   // assign rom_data[19029]=8'b00110111;
   // assign rom_data[19030]=8'b01000000;
   // assign rom_data[19031]=8'b00111001;
   // assign rom_data[19032]=8'b00111111;
   // assign rom_data[19033]=8'b00111010;
   // assign rom_data[19034]=8'b00111111;
   // assign rom_data[19035]=8'b00111011;
   // assign rom_data[19036]=8'b00111111;
   // assign rom_data[19037]=8'b00111100;
   // assign rom_data[19038]=8'b00111111;
   // assign rom_data[19039]=8'b00111101;
   // assign rom_data[19040]=8'b00111111;
   // assign rom_data[19041]=8'b00111110;
   // assign rom_data[19042]=8'b00111111;
   // assign rom_data[19043]=8'b01000000;
   // assign rom_data[19044]=8'b00111111;
   // assign rom_data[19045]=8'b01000001;
   // assign rom_data[19046]=8'b00111111;
   // assign rom_data[19047]=8'b01000010;
   // assign rom_data[19048]=8'b00111111;
   // assign rom_data[19049]=8'b01000100;
   // assign rom_data[19050]=8'b00111111;
   // assign rom_data[19051]=8'b01000101;
   // assign rom_data[19052]=8'b00111111;
   // assign rom_data[19053]=8'b01000110;
   // assign rom_data[19054]=8'b00111111;
   // assign rom_data[19055]=8'b01001000;
   // assign rom_data[19056]=8'b00111111;
   // assign rom_data[19057]=8'b01001001;
   // assign rom_data[19058]=8'b00111111;
   // assign rom_data[19059]=8'b01001010;
   // assign rom_data[19060]=8'b00111111;
   // assign rom_data[19061]=8'b01001100;
   // assign rom_data[19062]=8'b00111111;
   // assign rom_data[19063]=8'b01001101;
   // assign rom_data[19064]=8'b00111111;
   // assign rom_data[19065]=8'b01001110;
   // assign rom_data[19066]=8'b00111111;
   // assign rom_data[19067]=8'b01010000;
   // assign rom_data[19068]=8'b00111111;
   // assign rom_data[19069]=8'b01010001;
   // assign rom_data[19070]=8'b00111111;
   // assign rom_data[19071]=8'b01010011;
   // assign rom_data[19072]=8'b00111111;
   // assign rom_data[19073]=8'b01010100;
   // assign rom_data[19074]=8'b00111111;
   // assign rom_data[19075]=8'b01010101;
   // assign rom_data[19076]=8'b00111111;
   // assign rom_data[19077]=8'b01010111;
   // assign rom_data[19078]=8'b00111111;
   // assign rom_data[19079]=8'b01011000;
   // assign rom_data[19080]=8'b00111111;
   // assign rom_data[19081]=8'b01011010;
   // assign rom_data[19082]=8'b00111111;
   // assign rom_data[19083]=8'b01011011;
   // assign rom_data[19084]=8'b00111111;
   // assign rom_data[19085]=8'b01011100;
   // assign rom_data[19086]=8'b00111111;
   // assign rom_data[19087]=8'b01011110;
   // assign rom_data[19088]=8'b00111111;
   // assign rom_data[19089]=8'b01011111;
   // assign rom_data[19090]=8'b00111111;
   // assign rom_data[19091]=8'b01100001;
   // assign rom_data[19092]=8'b00111111;
   // assign rom_data[19093]=8'b01100010;
   // assign rom_data[19094]=8'b00111111;
   // assign rom_data[19095]=8'b01100011;
   // assign rom_data[19096]=8'b00111111;
   // assign rom_data[19097]=8'b01100101;
   // assign rom_data[19098]=8'b00111111;
   // assign rom_data[19099]=8'b01100110;
   // assign rom_data[19100]=8'b00111111;
   // assign rom_data[19101]=8'b01101000;
   // assign rom_data[19102]=8'b00111111;
   // assign rom_data[19103]=8'b01101001;
   // assign rom_data[19104]=8'b00111111;
   // assign rom_data[19105]=8'b01101010;
   // assign rom_data[19106]=8'b00111111;
   // assign rom_data[19107]=8'b01101100;
   // assign rom_data[19108]=8'b00111111;
   // assign rom_data[19109]=8'b01101101;
   // assign rom_data[19110]=8'b00111111;
   // assign rom_data[19111]=8'b01101110;
   // assign rom_data[19112]=8'b00111111;
   // assign rom_data[19113]=8'b01110000;
   // assign rom_data[19114]=8'b00111111;
   // assign rom_data[19115]=8'b01110001;
   // assign rom_data[19116]=8'b00111111;
   // assign rom_data[19117]=8'b01110010;
   // assign rom_data[19118]=8'b00111111;
   // assign rom_data[19119]=8'b01110100;
   // assign rom_data[19120]=8'b00111111;
   // assign rom_data[19121]=8'b01110101;
   // assign rom_data[19122]=8'b00111111;
   // assign rom_data[19123]=8'b01110110;
   // assign rom_data[19124]=8'b00111111;
   // assign rom_data[19125]=8'b01110111;
   // assign rom_data[19126]=8'b00111111;
   // assign rom_data[19127]=8'b01111001;
   // assign rom_data[19128]=8'b00111111;
   // assign rom_data[19129]=8'b01111010;
   // assign rom_data[19130]=8'b00111111;
   // assign rom_data[19131]=8'b01111011;
   // assign rom_data[19132]=8'b00111111;
   // assign rom_data[19133]=8'b01111100;
   // assign rom_data[19134]=8'b00111111;
   // assign rom_data[19135]=8'b01111101;
   // assign rom_data[19136]=8'b00111111;
   // assign rom_data[19137]=8'b01111110;
   // assign rom_data[19138]=8'b00111111;
   // assign rom_data[19139]=8'b01111111;
   // assign rom_data[19140]=8'b00111111;
   // assign rom_data[19141]=8'b10000000;
   // assign rom_data[19142]=8'b00111111;
   // assign rom_data[19143]=8'b10000001;
   // assign rom_data[19144]=8'b00111111;
   // assign rom_data[19145]=8'b10000010;
   // assign rom_data[19146]=8'b00111111;
   // assign rom_data[19147]=8'b10000011;
   // assign rom_data[19148]=8'b00111111;
   // assign rom_data[19149]=8'b10000100;
   // assign rom_data[19150]=8'b00111111;
   // assign rom_data[19151]=8'b10000101;
   // assign rom_data[19152]=8'b00111110;
   // assign rom_data[19153]=8'b10000110;
   // assign rom_data[19154]=8'b00111110;
   // assign rom_data[19155]=8'b10000110;
   // assign rom_data[19156]=8'b00111110;
   // assign rom_data[19157]=8'b10000111;
   // assign rom_data[19158]=8'b00111110;
   // assign rom_data[19159]=8'b10001000;
   // assign rom_data[19160]=8'b00111110;
   // assign rom_data[19161]=8'b10001000;
   // assign rom_data[19162]=8'b00111110;
   // assign rom_data[19163]=8'b10001001;
   // assign rom_data[19164]=8'b00111110;
   // assign rom_data[19165]=8'b10001001;
   // assign rom_data[19166]=8'b00111110;
   // assign rom_data[19167]=8'b10001001;
   // assign rom_data[19168]=8'b00111110;
   // assign rom_data[19169]=8'b10001010;
   // assign rom_data[19170]=8'b00111110;
   // assign rom_data[19171]=8'b10001010;
   // assign rom_data[19172]=8'b00111110;
   // assign rom_data[19173]=8'b10001010;
   // assign rom_data[19174]=8'b00111110;
   // assign rom_data[19175]=8'b10001010;
   // assign rom_data[19176]=8'b00111110;
   // assign rom_data[19177]=8'b10001010;
   // assign rom_data[19178]=8'b00111110;
   // assign rom_data[19179]=8'b10001001;
   // assign rom_data[19180]=8'b00111110;
   // assign rom_data[19181]=8'b10001001;
   // assign rom_data[19182]=8'b00111110;
   // assign rom_data[19183]=8'b10001001;
   // assign rom_data[19184]=8'b00111110;
   // assign rom_data[19185]=8'b10001000;
   // assign rom_data[19186]=8'b00111110;
   // assign rom_data[19187]=8'b10001000;
   // assign rom_data[19188]=8'b00111110;
   // assign rom_data[19189]=8'b10000111;
   // assign rom_data[19190]=8'b00111110;
   // assign rom_data[19191]=8'b10000111;
   // assign rom_data[19192]=8'b00111110;
   // assign rom_data[19193]=8'b10000110;
   // assign rom_data[19194]=8'b00111110;
   // assign rom_data[19195]=8'b10000101;
   // assign rom_data[19196]=8'b00111110;
   // assign rom_data[19197]=8'b10000100;
   // assign rom_data[19198]=8'b00111110;
   // assign rom_data[19199]=8'b10000011;
   // assign rom_data[19200]=8'b00111110;
   // assign rom_data[19201]=8'b10000010;
   // assign rom_data[19202]=8'b00111110;
   // assign rom_data[19203]=8'b10000010;
   // assign rom_data[19204]=8'b00111110;
   // assign rom_data[19205]=8'b10000001;
   // assign rom_data[19206]=8'b00111110;
   // assign rom_data[19207]=8'b01111111;
   // assign rom_data[19208]=8'b00111110;
   // assign rom_data[19209]=8'b01111110;
   // assign rom_data[19210]=8'b00111110;
   // assign rom_data[19211]=8'b01111101;
   // assign rom_data[19212]=8'b00111110;
   // assign rom_data[19213]=8'b01111100;
   // assign rom_data[19214]=8'b00111110;
   // assign rom_data[19215]=8'b01111011;
   // assign rom_data[19216]=8'b00111110;
   // assign rom_data[19217]=8'b01111010;
   // assign rom_data[19218]=8'b00111110;
   // assign rom_data[19219]=8'b01111001;
   // assign rom_data[19220]=8'b00111110;
   // assign rom_data[19221]=8'b01110111;
   // assign rom_data[19222]=8'b00111110;
   // assign rom_data[19223]=8'b01110110;
   // assign rom_data[19224]=8'b00111110;
   // assign rom_data[19225]=8'b01110101;
   // assign rom_data[19226]=8'b00111110;
   // assign rom_data[19227]=8'b01110100;
   // assign rom_data[19228]=8'b00111110;
   // assign rom_data[19229]=8'b01110010;
   // assign rom_data[19230]=8'b00111110;
   // assign rom_data[19231]=8'b01110001;
   // assign rom_data[19232]=8'b00111110;
   // assign rom_data[19233]=8'b01110000;
   // assign rom_data[19234]=8'b00111110;
   // assign rom_data[19235]=8'b01101110;
   // assign rom_data[19236]=8'b00111110;
   // assign rom_data[19237]=8'b01101101;
   // assign rom_data[19238]=8'b00111110;
   // assign rom_data[19239]=8'b01101100;
   // assign rom_data[19240]=8'b00111110;
   // assign rom_data[19241]=8'b01101010;
   // assign rom_data[19242]=8'b00111110;
   // assign rom_data[19243]=8'b01101001;
   // assign rom_data[19244]=8'b00111110;
   // assign rom_data[19245]=8'b01100111;
   // assign rom_data[19246]=8'b00111110;
   // assign rom_data[19247]=8'b01100110;
   // assign rom_data[19248]=8'b00111110;
   // assign rom_data[19249]=8'b01100101;
   // assign rom_data[19250]=8'b00111110;
   // assign rom_data[19251]=8'b01100011;
   // assign rom_data[19252]=8'b00111110;
   // assign rom_data[19253]=8'b01100010;
   // assign rom_data[19254]=8'b00111110;
   // assign rom_data[19255]=8'b01100000;
   // assign rom_data[19256]=8'b00111110;
   // assign rom_data[19257]=8'b01011111;
   // assign rom_data[19258]=8'b00111110;
   // assign rom_data[19259]=8'b01011110;
   // assign rom_data[19260]=8'b00111110;
   // assign rom_data[19261]=8'b01011100;
   // assign rom_data[19262]=8'b00111101;
   // assign rom_data[19263]=8'b01011011;
   // assign rom_data[19264]=8'b00111101;
   // assign rom_data[19265]=8'b01011001;
   // assign rom_data[19266]=8'b00111101;
   // assign rom_data[19267]=8'b01011000;
   // assign rom_data[19268]=8'b00111101;
   // assign rom_data[19269]=8'b01010111;
   // assign rom_data[19270]=8'b00111101;
   // assign rom_data[19271]=8'b01010101;
   // assign rom_data[19272]=8'b00111101;
   // assign rom_data[19273]=8'b01010100;
   // assign rom_data[19274]=8'b00111101;
   // assign rom_data[19275]=8'b01010010;
   // assign rom_data[19276]=8'b00111101;
   // assign rom_data[19277]=8'b01010001;
   // assign rom_data[19278]=8'b00111101;
   // assign rom_data[19279]=8'b01010000;
   // assign rom_data[19280]=8'b00111101;
   // assign rom_data[19281]=8'b01001110;
   // assign rom_data[19282]=8'b00111101;
   // assign rom_data[19283]=8'b01001101;
   // assign rom_data[19284]=8'b00111101;
   // assign rom_data[19285]=8'b01001100;
   // assign rom_data[19286]=8'b00111101;
   // assign rom_data[19287]=8'b01001010;
   // assign rom_data[19288]=8'b00111101;
   // assign rom_data[19289]=8'b01001001;
   // assign rom_data[19290]=8'b00111101;
   // assign rom_data[19291]=8'b01000111;
   // assign rom_data[19292]=8'b00111101;
   // assign rom_data[19293]=8'b01000110;
   // assign rom_data[19294]=8'b00111101;
   // assign rom_data[19295]=8'b01000101;
   // assign rom_data[19296]=8'b00111101;
   // assign rom_data[19297]=8'b01000100;
   // assign rom_data[19298]=8'b00111101;
   // assign rom_data[19299]=8'b01000010;
   // assign rom_data[19300]=8'b00111101;
   // assign rom_data[19301]=8'b01000001;
   // assign rom_data[19302]=8'b00111101;
   // assign rom_data[19303]=8'b01000000;
   // assign rom_data[19304]=8'b00111101;
   // assign rom_data[19305]=8'b00111110;
   // assign rom_data[19306]=8'b00111101;
   // assign rom_data[19307]=8'b00111101;
   // assign rom_data[19308]=8'b00111101;
   // assign rom_data[19309]=8'b00111100;
   // assign rom_data[19310]=8'b00111101;
   // assign rom_data[19311]=8'b00111011;
   // assign rom_data[19312]=8'b00111101;
   // assign rom_data[19313]=8'b00111010;
   // assign rom_data[19314]=8'b00111101;
   // assign rom_data[19315]=8'b00111001;
   // assign rom_data[19316]=8'b00111101;
   // assign rom_data[19317]=8'b00110111;
   // assign rom_data[19318]=8'b00111101;
   // assign rom_data[19319]=8'b00110110;
   // assign rom_data[19320]=8'b00111101;
   // assign rom_data[19321]=8'b00110101;
   // assign rom_data[19322]=8'b00111101;
   // assign rom_data[19323]=8'b00110100;
   // assign rom_data[19324]=8'b00111101;
   // assign rom_data[19325]=8'b00110011;
   // assign rom_data[19326]=8'b00111101;
   // assign rom_data[19327]=8'b00110010;
   // assign rom_data[19328]=8'b00111101;
   // assign rom_data[19329]=8'b00110010;
   // assign rom_data[19330]=8'b00111101;
   // assign rom_data[19331]=8'b00110001;
   // assign rom_data[19332]=8'b00111101;
   // assign rom_data[19333]=8'b00110000;
   // assign rom_data[19334]=8'b00111101;
   // assign rom_data[19335]=8'b00101111;
   // assign rom_data[19336]=8'b00111101;
   // assign rom_data[19337]=8'b00101111;
   // assign rom_data[19338]=8'b00111101;
   // assign rom_data[19339]=8'b00101110;
   // assign rom_data[19340]=8'b00111101;
   // assign rom_data[19341]=8'b00101110;
   // assign rom_data[19342]=8'b00111101;
   // assign rom_data[19343]=8'b00101101;
   // assign rom_data[19344]=8'b00111101;
   // assign rom_data[19345]=8'b00101101;
   // assign rom_data[19346]=8'b00111101;
   // assign rom_data[19347]=8'b00101100;
   // assign rom_data[19348]=8'b00111101;
   // assign rom_data[19349]=8'b00101100;
   // assign rom_data[19350]=8'b00111101;
   // assign rom_data[19351]=8'b00101100;
   // assign rom_data[19352]=8'b00111101;
   // assign rom_data[19353]=8'b00101100;
   // assign rom_data[19354]=8'b00111101;
   // assign rom_data[19355]=8'b00101100;
   // assign rom_data[19356]=8'b00111101;
   // assign rom_data[19357]=8'b00101100;
   // assign rom_data[19358]=8'b00111101;
   // assign rom_data[19359]=8'b00101100;
   // assign rom_data[19360]=8'b00111101;
   // assign rom_data[19361]=8'b00101101;
   // assign rom_data[19362]=8'b00111101;
   // assign rom_data[19363]=8'b00101101;
   // assign rom_data[19364]=8'b00111101;
   // assign rom_data[19365]=8'b00101101;
   // assign rom_data[19366]=8'b00111101;
   // assign rom_data[19367]=8'b00101110;
   // assign rom_data[19368]=8'b00111101;
   // assign rom_data[19369]=8'b00101111;
   // assign rom_data[19370]=8'b00111101;
   // assign rom_data[19371]=8'b00101111;
   // assign rom_data[19372]=8'b00111100;
   // assign rom_data[19373]=8'b00110000;
   // assign rom_data[19374]=8'b00111100;
   // assign rom_data[19375]=8'b00110001;
   // assign rom_data[19376]=8'b00111100;
   // assign rom_data[19377]=8'b00110010;
   // assign rom_data[19378]=8'b00111100;
   // assign rom_data[19379]=8'b00110010;
   // assign rom_data[19380]=8'b00111100;
   // assign rom_data[19381]=8'b00110011;
   // assign rom_data[19382]=8'b00111100;
   // assign rom_data[19383]=8'b00110100;
   // assign rom_data[19384]=8'b00111100;
   // assign rom_data[19385]=8'b00110101;
   // assign rom_data[19386]=8'b00111100;
   // assign rom_data[19387]=8'b00110110;
   // assign rom_data[19388]=8'b00111100;
   // assign rom_data[19389]=8'b00110111;
   // assign rom_data[19390]=8'b00111100;
   // assign rom_data[19391]=8'b00111001;
   // assign rom_data[19392]=8'b00111100;
   // assign rom_data[19393]=8'b00111010;
   // assign rom_data[19394]=8'b00111100;
   // assign rom_data[19395]=8'b00111011;
   // assign rom_data[19396]=8'b00111100;
   // assign rom_data[19397]=8'b00111100;
   // assign rom_data[19398]=8'b00111100;
   // assign rom_data[19399]=8'b00111101;
   // assign rom_data[19400]=8'b00111100;
   // assign rom_data[19401]=8'b00111110;
   // assign rom_data[19402]=8'b00111100;
   // assign rom_data[19403]=8'b01000000;
   // assign rom_data[19404]=8'b00111100;
   // assign rom_data[19405]=8'b01000001;
   // assign rom_data[19406]=8'b00111100;
   // assign rom_data[19407]=8'b01000010;
   // assign rom_data[19408]=8'b00111100;
   // assign rom_data[19409]=8'b01000100;
   // assign rom_data[19410]=8'b00111100;
   // assign rom_data[19411]=8'b01000101;
   // assign rom_data[19412]=8'b00111100;
   // assign rom_data[19413]=8'b01000110;
   // assign rom_data[19414]=8'b00111100;
   // assign rom_data[19415]=8'b01001000;
   // assign rom_data[19416]=8'b00111100;
   // assign rom_data[19417]=8'b01001001;
   // assign rom_data[19418]=8'b00111100;
   // assign rom_data[19419]=8'b01001010;
   // assign rom_data[19420]=8'b00111100;
   // assign rom_data[19421]=8'b01001100;
   // assign rom_data[19422]=8'b00111100;
   // assign rom_data[19423]=8'b01001101;
   // assign rom_data[19424]=8'b00111100;
   // assign rom_data[19425]=8'b01001110;
   // assign rom_data[19426]=8'b00111100;
   // assign rom_data[19427]=8'b01010000;
   // assign rom_data[19428]=8'b00111100;
   // assign rom_data[19429]=8'b01010001;
   // assign rom_data[19430]=8'b00111100;
   // assign rom_data[19431]=8'b01010011;
   // assign rom_data[19432]=8'b00111100;
   // assign rom_data[19433]=8'b01010100;
   // assign rom_data[19434]=8'b00111100;
   // assign rom_data[19435]=8'b01010101;
   // assign rom_data[19436]=8'b00111100;
   // assign rom_data[19437]=8'b01010111;
   // assign rom_data[19438]=8'b00111100;
   // assign rom_data[19439]=8'b01011000;
   // assign rom_data[19440]=8'b00111100;
   // assign rom_data[19441]=8'b01011010;
   // assign rom_data[19442]=8'b00111100;
   // assign rom_data[19443]=8'b01011011;
   // assign rom_data[19444]=8'b00111100;
   // assign rom_data[19445]=8'b01011100;
   // assign rom_data[19446]=8'b00111100;
   // assign rom_data[19447]=8'b01011110;
   // assign rom_data[19448]=8'b00111100;
   // assign rom_data[19449]=8'b01011111;
   // assign rom_data[19450]=8'b00111100;
   // assign rom_data[19451]=8'b01100001;
   // assign rom_data[19452]=8'b00111100;
   // assign rom_data[19453]=8'b01100010;
   // assign rom_data[19454]=8'b00111100;
   // assign rom_data[19455]=8'b01100011;
   // assign rom_data[19456]=8'b00111100;
   // assign rom_data[19457]=8'b01100101;
   // assign rom_data[19458]=8'b00111100;
   // assign rom_data[19459]=8'b01100110;
   // assign rom_data[19460]=8'b00111100;
   // assign rom_data[19461]=8'b01101000;
   // assign rom_data[19462]=8'b00111100;
   // assign rom_data[19463]=8'b01101001;
   // assign rom_data[19464]=8'b00111100;
   // assign rom_data[19465]=8'b01101010;
   // assign rom_data[19466]=8'b00111100;
   // assign rom_data[19467]=8'b01101100;
   // assign rom_data[19468]=8'b00111100;
   // assign rom_data[19469]=8'b01101101;
   // assign rom_data[19470]=8'b00111100;
   // assign rom_data[19471]=8'b01101110;
   // assign rom_data[19472]=8'b00111100;
   // assign rom_data[19473]=8'b01110000;
   // assign rom_data[19474]=8'b00111100;
   // assign rom_data[19475]=8'b01110001;
   // assign rom_data[19476]=8'b00111100;
   // assign rom_data[19477]=8'b01110010;
   // assign rom_data[19478]=8'b00111100;
   // assign rom_data[19479]=8'b01110100;
   // assign rom_data[19480]=8'b00111100;
   // assign rom_data[19481]=8'b01110101;
   // assign rom_data[19482]=8'b00111100;
   // assign rom_data[19483]=8'b01110110;
   // assign rom_data[19484]=8'b00111100;
   // assign rom_data[19485]=8'b01110111;
   // assign rom_data[19486]=8'b00111100;
   // assign rom_data[19487]=8'b01111001;
   // assign rom_data[19488]=8'b00111100;
   // assign rom_data[19489]=8'b01111010;
   // assign rom_data[19490]=8'b00111100;
   // assign rom_data[19491]=8'b01111011;
   // assign rom_data[19492]=8'b00111100;
   // assign rom_data[19493]=8'b01111100;
   // assign rom_data[19494]=8'b00111011;
   // assign rom_data[19495]=8'b01111101;
   // assign rom_data[19496]=8'b00111011;
   // assign rom_data[19497]=8'b01111110;
   // assign rom_data[19498]=8'b00111011;
   // assign rom_data[19499]=8'b01111111;
   // assign rom_data[19500]=8'b00111011;
   // assign rom_data[19501]=8'b10000000;
   // assign rom_data[19502]=8'b00111011;
   // assign rom_data[19503]=8'b10000001;
   // assign rom_data[19504]=8'b00111011;
   // assign rom_data[19505]=8'b10000010;
   // assign rom_data[19506]=8'b00111011;
   // assign rom_data[19507]=8'b10000011;
   // assign rom_data[19508]=8'b00111011;
   // assign rom_data[19509]=8'b10000100;
   // assign rom_data[19510]=8'b00111011;
   // assign rom_data[19511]=8'b10000101;
   // assign rom_data[19512]=8'b00111011;
   // assign rom_data[19513]=8'b10000110;
   // assign rom_data[19514]=8'b00111011;
   // assign rom_data[19515]=8'b10000110;
   // assign rom_data[19516]=8'b00111011;
   // assign rom_data[19517]=8'b10000111;
   // assign rom_data[19518]=8'b00111011;
   // assign rom_data[19519]=8'b10001000;
   // assign rom_data[19520]=8'b00111011;
   // assign rom_data[19521]=8'b10001000;
   // assign rom_data[19522]=8'b00111011;
   // assign rom_data[19523]=8'b10001001;
   // assign rom_data[19524]=8'b00111011;
   // assign rom_data[19525]=8'b10001001;
   // assign rom_data[19526]=8'b00111011;
   // assign rom_data[19527]=8'b10001001;
   // assign rom_data[19528]=8'b00111011;
   // assign rom_data[19529]=8'b10001010;
   // assign rom_data[19530]=8'b00111011;
   // assign rom_data[19531]=8'b10001010;
   // assign rom_data[19532]=8'b00111011;
   // assign rom_data[19533]=8'b10001010;
   // assign rom_data[19534]=8'b00111011;
   // assign rom_data[19535]=8'b10001010;
   // assign rom_data[19536]=8'b00111011;
   // assign rom_data[19537]=8'b10001010;
   // assign rom_data[19538]=8'b00111011;
   // assign rom_data[19539]=8'b10001001;
   // assign rom_data[19540]=8'b00111011;
   // assign rom_data[19541]=8'b10001001;
   // assign rom_data[19542]=8'b00111011;
   // assign rom_data[19543]=8'b10001001;
   // assign rom_data[19544]=8'b00111011;
   // assign rom_data[19545]=8'b10001000;
   // assign rom_data[19546]=8'b00111011;
   // assign rom_data[19547]=8'b10001000;
   // assign rom_data[19548]=8'b00111011;
   // assign rom_data[19549]=8'b10000111;
   // assign rom_data[19550]=8'b00111011;
   // assign rom_data[19551]=8'b10000111;
   // assign rom_data[19552]=8'b00111011;
   // assign rom_data[19553]=8'b10000110;
   // assign rom_data[19554]=8'b00111011;
   // assign rom_data[19555]=8'b10000101;
   // assign rom_data[19556]=8'b00111011;
   // assign rom_data[19557]=8'b10000100;
   // assign rom_data[19558]=8'b00111011;
   // assign rom_data[19559]=8'b10000011;
   // assign rom_data[19560]=8'b00111011;
   // assign rom_data[19561]=8'b10000010;
   // assign rom_data[19562]=8'b00111011;
   // assign rom_data[19563]=8'b10000010;
   // assign rom_data[19564]=8'b00111011;
   // assign rom_data[19565]=8'b10000001;
   // assign rom_data[19566]=8'b00111011;
   // assign rom_data[19567]=8'b01111111;
   // assign rom_data[19568]=8'b00111011;
   // assign rom_data[19569]=8'b01111110;
   // assign rom_data[19570]=8'b00111011;
   // assign rom_data[19571]=8'b01111101;
   // assign rom_data[19572]=8'b00111011;
   // assign rom_data[19573]=8'b01111100;
   // assign rom_data[19574]=8'b00111011;
   // assign rom_data[19575]=8'b01111011;
   // assign rom_data[19576]=8'b00111011;
   // assign rom_data[19577]=8'b01111010;
   // assign rom_data[19578]=8'b00111011;
   // assign rom_data[19579]=8'b01111001;
   // assign rom_data[19580]=8'b00111011;
   // assign rom_data[19581]=8'b01110111;
   // assign rom_data[19582]=8'b00111011;
   // assign rom_data[19583]=8'b01110110;
   // assign rom_data[19584]=8'b00111011;
   // assign rom_data[19585]=8'b01110101;
   // assign rom_data[19586]=8'b00111011;
   // assign rom_data[19587]=8'b01110100;
   // assign rom_data[19588]=8'b00111011;
   // assign rom_data[19589]=8'b01110010;
   // assign rom_data[19590]=8'b00111011;
   // assign rom_data[19591]=8'b01110001;
   // assign rom_data[19592]=8'b00111011;
   // assign rom_data[19593]=8'b01110000;
   // assign rom_data[19594]=8'b00111011;
   // assign rom_data[19595]=8'b01101110;
   // assign rom_data[19596]=8'b00111011;
   // assign rom_data[19597]=8'b01101101;
   // assign rom_data[19598]=8'b00111011;
   // assign rom_data[19599]=8'b01101100;
   // assign rom_data[19600]=8'b00111010;
   // assign rom_data[19601]=8'b01101010;
   // assign rom_data[19602]=8'b00111010;
   // assign rom_data[19603]=8'b01101001;
   // assign rom_data[19604]=8'b00111010;
   // assign rom_data[19605]=8'b01100111;
   // assign rom_data[19606]=8'b00111010;
   // assign rom_data[19607]=8'b01100110;
   // assign rom_data[19608]=8'b00111010;
   // assign rom_data[19609]=8'b01100101;
   // assign rom_data[19610]=8'b00111010;
   // assign rom_data[19611]=8'b01100011;
   // assign rom_data[19612]=8'b00111010;
   // assign rom_data[19613]=8'b01100010;
   // assign rom_data[19614]=8'b00111010;
   // assign rom_data[19615]=8'b01100000;
   // assign rom_data[19616]=8'b00111010;
   // assign rom_data[19617]=8'b01011111;
   // assign rom_data[19618]=8'b00111010;
   // assign rom_data[19619]=8'b01011110;
   // assign rom_data[19620]=8'b00111010;
   // assign rom_data[19621]=8'b01011100;
   // assign rom_data[19622]=8'b00111010;
   // assign rom_data[19623]=8'b01011011;
   // assign rom_data[19624]=8'b00111010;
   // assign rom_data[19625]=8'b01011001;
   // assign rom_data[19626]=8'b00111010;
   // assign rom_data[19627]=8'b01011000;
   // assign rom_data[19628]=8'b00111010;
   // assign rom_data[19629]=8'b01010111;
   // assign rom_data[19630]=8'b00111010;
   // assign rom_data[19631]=8'b01010101;
   // assign rom_data[19632]=8'b00111010;
   // assign rom_data[19633]=8'b01010100;
   // assign rom_data[19634]=8'b00111010;
   // assign rom_data[19635]=8'b01010010;
   // assign rom_data[19636]=8'b00111010;
   // assign rom_data[19637]=8'b01010001;
   // assign rom_data[19638]=8'b00111010;
   // assign rom_data[19639]=8'b01010000;
   // assign rom_data[19640]=8'b00111010;
   // assign rom_data[19641]=8'b01001110;
   // assign rom_data[19642]=8'b00111010;
   // assign rom_data[19643]=8'b01001101;
   // assign rom_data[19644]=8'b00111010;
   // assign rom_data[19645]=8'b01001100;
   // assign rom_data[19646]=8'b00111010;
   // assign rom_data[19647]=8'b01001010;
   // assign rom_data[19648]=8'b00111010;
   // assign rom_data[19649]=8'b01001001;
   // assign rom_data[19650]=8'b00111010;
   // assign rom_data[19651]=8'b01000111;
   // assign rom_data[19652]=8'b00111010;
   // assign rom_data[19653]=8'b01000110;
   // assign rom_data[19654]=8'b00111010;
   // assign rom_data[19655]=8'b01000101;
   // assign rom_data[19656]=8'b00111010;
   // assign rom_data[19657]=8'b01000100;
   // assign rom_data[19658]=8'b00111010;
   // assign rom_data[19659]=8'b01000010;
   // assign rom_data[19660]=8'b00111010;
   // assign rom_data[19661]=8'b01000001;
   // assign rom_data[19662]=8'b00111010;
   // assign rom_data[19663]=8'b01000000;
   // assign rom_data[19664]=8'b00111010;
   // assign rom_data[19665]=8'b00111110;
   // assign rom_data[19666]=8'b00111010;
   // assign rom_data[19667]=8'b00111101;
   // assign rom_data[19668]=8'b00111010;
   // assign rom_data[19669]=8'b00111100;
   // assign rom_data[19670]=8'b00111010;
   // assign rom_data[19671]=8'b00111011;
   // assign rom_data[19672]=8'b00111010;
   // assign rom_data[19673]=8'b00111010;
   // assign rom_data[19674]=8'b00111010;
   // assign rom_data[19675]=8'b00111001;
   // assign rom_data[19676]=8'b00111010;
   // assign rom_data[19677]=8'b00110111;
   // assign rom_data[19678]=8'b00111010;
   // assign rom_data[19679]=8'b00110110;
   // assign rom_data[19680]=8'b00111010;
   // assign rom_data[19681]=8'b00110101;
   // assign rom_data[19682]=8'b00111010;
   // assign rom_data[19683]=8'b00110100;
   // assign rom_data[19684]=8'b00111010;
   // assign rom_data[19685]=8'b00110011;
   // assign rom_data[19686]=8'b00111010;
   // assign rom_data[19687]=8'b00110010;
   // assign rom_data[19688]=8'b00111010;
   // assign rom_data[19689]=8'b00110010;
   // assign rom_data[19690]=8'b00111010;
   // assign rom_data[19691]=8'b00110001;
   // assign rom_data[19692]=8'b00111010;
   // assign rom_data[19693]=8'b00110000;
   // assign rom_data[19694]=8'b00111010;
   // assign rom_data[19695]=8'b00101111;
   // assign rom_data[19696]=8'b00111010;
   // assign rom_data[19697]=8'b00101111;
   // assign rom_data[19698]=8'b00111010;
   // assign rom_data[19699]=8'b00101110;
   // assign rom_data[19700]=8'b00111010;
   // assign rom_data[19701]=8'b00101110;
   // assign rom_data[19702]=8'b00111010;
   // assign rom_data[19703]=8'b00101101;
   // assign rom_data[19704]=8'b00111010;
   // assign rom_data[19705]=8'b00101101;
   // assign rom_data[19706]=8'b00111010;
   // assign rom_data[19707]=8'b00101100;
   // assign rom_data[19708]=8'b00111010;
   // assign rom_data[19709]=8'b00101100;
   // assign rom_data[19710]=8'b00111010;
   // assign rom_data[19711]=8'b00101100;
   // assign rom_data[19712]=8'b00111010;
   // assign rom_data[19713]=8'b00101100;
   // assign rom_data[19714]=8'b00111001;
   // assign rom_data[19715]=8'b00101100;
   // assign rom_data[19716]=8'b00111001;
   // assign rom_data[19717]=8'b00101100;
   // assign rom_data[19718]=8'b00111001;
   // assign rom_data[19719]=8'b00101100;
   // assign rom_data[19720]=8'b00111001;
   // assign rom_data[19721]=8'b00101101;
   // assign rom_data[19722]=8'b00111001;
   // assign rom_data[19723]=8'b00101101;
   // assign rom_data[19724]=8'b00111001;
   // assign rom_data[19725]=8'b00101101;
   // assign rom_data[19726]=8'b00111001;
   // assign rom_data[19727]=8'b00101110;
   // assign rom_data[19728]=8'b00111001;
   // assign rom_data[19729]=8'b00101111;
   // assign rom_data[19730]=8'b00111001;
   // assign rom_data[19731]=8'b00101111;
   // assign rom_data[19732]=8'b00111001;
   // assign rom_data[19733]=8'b00110000;
   // assign rom_data[19734]=8'b00111001;
   // assign rom_data[19735]=8'b00110001;
   // assign rom_data[19736]=8'b00111001;
   // assign rom_data[19737]=8'b00110010;
   // assign rom_data[19738]=8'b00111001;
   // assign rom_data[19739]=8'b00110010;
   // assign rom_data[19740]=8'b00111001;
   // assign rom_data[19741]=8'b00110011;
   // assign rom_data[19742]=8'b00111001;
   // assign rom_data[19743]=8'b00110100;
   // assign rom_data[19744]=8'b00111001;
   // assign rom_data[19745]=8'b00110101;
   // assign rom_data[19746]=8'b00111001;
   // assign rom_data[19747]=8'b00110110;
   // assign rom_data[19748]=8'b00111001;
   // assign rom_data[19749]=8'b00110111;
   // assign rom_data[19750]=8'b00111001;
   // assign rom_data[19751]=8'b00111001;
   // assign rom_data[19752]=8'b00111001;
   // assign rom_data[19753]=8'b00111010;
   // assign rom_data[19754]=8'b00111001;
   // assign rom_data[19755]=8'b00111011;
   // assign rom_data[19756]=8'b00111001;
   // assign rom_data[19757]=8'b00111100;
   // assign rom_data[19758]=8'b00111001;
   // assign rom_data[19759]=8'b00111101;
   // assign rom_data[19760]=8'b00111001;
   // assign rom_data[19761]=8'b00111110;
   // assign rom_data[19762]=8'b00111001;
   // assign rom_data[19763]=8'b01000000;
   // assign rom_data[19764]=8'b00111001;
   // assign rom_data[19765]=8'b01000001;
   // assign rom_data[19766]=8'b00111001;
   // assign rom_data[19767]=8'b01000010;
   // assign rom_data[19768]=8'b00111001;
   // assign rom_data[19769]=8'b01000100;
   // assign rom_data[19770]=8'b00111001;
   // assign rom_data[19771]=8'b01000101;
   // assign rom_data[19772]=8'b00111001;
   // assign rom_data[19773]=8'b01000110;
   // assign rom_data[19774]=8'b00111001;
   // assign rom_data[19775]=8'b01001000;
   // assign rom_data[19776]=8'b00111001;
   // assign rom_data[19777]=8'b01001001;
   // assign rom_data[19778]=8'b00111001;
   // assign rom_data[19779]=8'b01001010;
   // assign rom_data[19780]=8'b00111001;
   // assign rom_data[19781]=8'b01001100;
   // assign rom_data[19782]=8'b00111001;
   // assign rom_data[19783]=8'b01001101;
   // assign rom_data[19784]=8'b00111001;
   // assign rom_data[19785]=8'b01001110;
   // assign rom_data[19786]=8'b00111001;
   // assign rom_data[19787]=8'b01010000;
   // assign rom_data[19788]=8'b00111001;
   // assign rom_data[19789]=8'b01010001;
   // assign rom_data[19790]=8'b00111001;
   // assign rom_data[19791]=8'b01010011;
   // assign rom_data[19792]=8'b00111001;
   // assign rom_data[19793]=8'b01010100;
   // assign rom_data[19794]=8'b00111001;
   // assign rom_data[19795]=8'b01010101;
   // assign rom_data[19796]=8'b00111001;
   // assign rom_data[19797]=8'b01010111;
   // assign rom_data[19798]=8'b00111001;
   // assign rom_data[19799]=8'b01011000;
   // assign rom_data[19800]=8'b00111001;
   // assign rom_data[19801]=8'b01011010;
   // assign rom_data[19802]=8'b00111001;
   // assign rom_data[19803]=8'b01011011;
   // assign rom_data[19804]=8'b00111001;
   // assign rom_data[19805]=8'b01011100;
   // assign rom_data[19806]=8'b00111001;
   // assign rom_data[19807]=8'b01011110;
   // assign rom_data[19808]=8'b00111001;
   // assign rom_data[19809]=8'b01011111;
   // assign rom_data[19810]=8'b00111001;
   // assign rom_data[19811]=8'b01100001;
   // assign rom_data[19812]=8'b00111001;
   // assign rom_data[19813]=8'b01100010;
   // assign rom_data[19814]=8'b00111001;
   // assign rom_data[19815]=8'b01100011;
   // assign rom_data[19816]=8'b00111001;
   // assign rom_data[19817]=8'b01100101;
   // assign rom_data[19818]=8'b00111001;
   // assign rom_data[19819]=8'b01100110;
   // assign rom_data[19820]=8'b00111001;
   // assign rom_data[19821]=8'b01101000;
   // assign rom_data[19822]=8'b00111001;
   // assign rom_data[19823]=8'b01101001;
   // assign rom_data[19824]=8'b00111001;
   // assign rom_data[19825]=8'b01101010;
   // assign rom_data[19826]=8'b00111001;
   // assign rom_data[19827]=8'b01101100;
   // assign rom_data[19828]=8'b00111001;
   // assign rom_data[19829]=8'b01101101;
   // assign rom_data[19830]=8'b00111001;
   // assign rom_data[19831]=8'b01101110;
   // assign rom_data[19832]=8'b00111000;
   // assign rom_data[19833]=8'b01110000;
   // assign rom_data[19834]=8'b00111000;
   // assign rom_data[19835]=8'b01110001;
   // assign rom_data[19836]=8'b00111000;
   // assign rom_data[19837]=8'b01110010;
   // assign rom_data[19838]=8'b00111000;
   // assign rom_data[19839]=8'b01110100;
   // assign rom_data[19840]=8'b00111000;
   // assign rom_data[19841]=8'b01110101;
   // assign rom_data[19842]=8'b00111000;
   // assign rom_data[19843]=8'b01110110;
   // assign rom_data[19844]=8'b00111000;
   // assign rom_data[19845]=8'b01110111;
   // assign rom_data[19846]=8'b00111000;
   // assign rom_data[19847]=8'b01111001;
   // assign rom_data[19848]=8'b00111000;
   // assign rom_data[19849]=8'b01111010;
   // assign rom_data[19850]=8'b00111000;
   // assign rom_data[19851]=8'b01111011;
   // assign rom_data[19852]=8'b00111000;
   // assign rom_data[19853]=8'b01111100;
   // assign rom_data[19854]=8'b00111000;
   // assign rom_data[19855]=8'b01111101;
   // assign rom_data[19856]=8'b00111000;
   // assign rom_data[19857]=8'b01111110;
   // assign rom_data[19858]=8'b00111000;
   // assign rom_data[19859]=8'b01111111;
   // assign rom_data[19860]=8'b00111000;
   // assign rom_data[19861]=8'b10000000;
   // assign rom_data[19862]=8'b00111000;
   // assign rom_data[19863]=8'b10000001;
   // assign rom_data[19864]=8'b00111000;
   // assign rom_data[19865]=8'b10000010;
   // assign rom_data[19866]=8'b00111000;
   // assign rom_data[19867]=8'b10000011;
   // assign rom_data[19868]=8'b00111000;
   // assign rom_data[19869]=8'b10000100;
   // assign rom_data[19870]=8'b00111000;
   // assign rom_data[19871]=8'b10000101;
   // assign rom_data[19872]=8'b00111000;
   // assign rom_data[19873]=8'b10000110;
   // assign rom_data[19874]=8'b00111000;
   // assign rom_data[19875]=8'b10000110;
   // assign rom_data[19876]=8'b00111000;
   // assign rom_data[19877]=8'b10000111;
   // assign rom_data[19878]=8'b00111000;
   // assign rom_data[19879]=8'b10001000;
   // assign rom_data[19880]=8'b00111000;
   // assign rom_data[19881]=8'b10001000;
   // assign rom_data[19882]=8'b00111000;
   // assign rom_data[19883]=8'b10001001;
   // assign rom_data[19884]=8'b00111000;
   // assign rom_data[19885]=8'b10001001;
   // assign rom_data[19886]=8'b00111000;
   // assign rom_data[19887]=8'b10001001;
   // assign rom_data[19888]=8'b00111000;
   // assign rom_data[19889]=8'b10001010;
   // assign rom_data[19890]=8'b00111000;
   // assign rom_data[19891]=8'b10001010;
   // assign rom_data[19892]=8'b00111000;
   // assign rom_data[19893]=8'b10001010;
   // assign rom_data[19894]=8'b00111000;
   // assign rom_data[19895]=8'b10001010;
   // assign rom_data[19896]=8'b00111000;
   // assign rom_data[19897]=8'b10001010;
   // assign rom_data[19898]=8'b00111000;
   // assign rom_data[19899]=8'b10001001;
   // assign rom_data[19900]=8'b00111000;
   // assign rom_data[19901]=8'b10001001;
   // assign rom_data[19902]=8'b00111000;
   // assign rom_data[19903]=8'b10001001;
   // assign rom_data[19904]=8'b00111000;
   // assign rom_data[19905]=8'b10001000;
   // assign rom_data[19906]=8'b00111000;
   // assign rom_data[19907]=8'b10001000;
   // assign rom_data[19908]=8'b00111000;
   // assign rom_data[19909]=8'b10000111;
   // assign rom_data[19910]=8'b00111000;
   // assign rom_data[19911]=8'b10000111;
   // assign rom_data[19912]=8'b00111000;
   // assign rom_data[19913]=8'b10000110;
   // assign rom_data[19914]=8'b00111000;
   // assign rom_data[19915]=8'b10000101;
   // assign rom_data[19916]=8'b00111000;
   // assign rom_data[19917]=8'b10000100;
   // assign rom_data[19918]=8'b00111000;
   // assign rom_data[19919]=8'b10000011;
   // assign rom_data[19920]=8'b00111000;
   // assign rom_data[19921]=8'b10000010;
   // assign rom_data[19922]=8'b00111000;
   // assign rom_data[19923]=8'b10000010;
   // assign rom_data[19924]=8'b00111000;
   // assign rom_data[19925]=8'b10000001;
   // assign rom_data[19926]=8'b00111000;
   // assign rom_data[19927]=8'b01111111;
   // assign rom_data[19928]=8'b00111000;
   // assign rom_data[19929]=8'b01111110;
   // assign rom_data[19930]=8'b00111000;
   // assign rom_data[19931]=8'b01111101;
   // assign rom_data[19932]=8'b00111000;
   // assign rom_data[19933]=8'b01111100;
   // assign rom_data[19934]=8'b00111000;
   // assign rom_data[19935]=8'b01111011;
   // assign rom_data[19936]=8'b00111000;
   // assign rom_data[19937]=8'b01111010;
   // assign rom_data[19938]=8'b00110111;
   // assign rom_data[19939]=8'b01111001;
   // assign rom_data[19940]=8'b00110111;
   // assign rom_data[19941]=8'b01110111;
   // assign rom_data[19942]=8'b00110111;
   // assign rom_data[19943]=8'b01110110;
   // assign rom_data[19944]=8'b00110111;
   // assign rom_data[19945]=8'b01110101;
   // assign rom_data[19946]=8'b00110111;
   // assign rom_data[19947]=8'b01110100;
   // assign rom_data[19948]=8'b00110111;
   // assign rom_data[19949]=8'b01110010;
   // assign rom_data[19950]=8'b00110111;
   // assign rom_data[19951]=8'b01110001;
   // assign rom_data[19952]=8'b00110111;
   // assign rom_data[19953]=8'b01110000;
   // assign rom_data[19954]=8'b00110111;
   // assign rom_data[19955]=8'b01101110;
   // assign rom_data[19956]=8'b00110111;
   // assign rom_data[19957]=8'b01101101;
   // assign rom_data[19958]=8'b00110111;
   // assign rom_data[19959]=8'b01101100;
   // assign rom_data[19960]=8'b00110111;
   // assign rom_data[19961]=8'b01101010;
   // assign rom_data[19962]=8'b00110111;
   // assign rom_data[19963]=8'b01101001;
   // assign rom_data[19964]=8'b00110111;
   // assign rom_data[19965]=8'b01100111;
   // assign rom_data[19966]=8'b00110111;
   // assign rom_data[19967]=8'b01100110;
   // assign rom_data[19968]=8'b00110111;
   // assign rom_data[19969]=8'b01100101;
   // assign rom_data[19970]=8'b00110111;
   // assign rom_data[19971]=8'b01100011;
   // assign rom_data[19972]=8'b00110111;
   // assign rom_data[19973]=8'b01100010;
   // assign rom_data[19974]=8'b00110111;
   // assign rom_data[19975]=8'b01100000;
   // assign rom_data[19976]=8'b00110111;
   // assign rom_data[19977]=8'b01011111;
   // assign rom_data[19978]=8'b00110111;
   // assign rom_data[19979]=8'b01011110;
   // assign rom_data[19980]=8'b00110111;
   // assign rom_data[19981]=8'b01011100;
   // assign rom_data[19982]=8'b00110111;
   // assign rom_data[19983]=8'b01011011;
   // assign rom_data[19984]=8'b00110111;
   // assign rom_data[19985]=8'b01011001;
   // assign rom_data[19986]=8'b00110111;
   // assign rom_data[19987]=8'b01011000;
   // assign rom_data[19988]=8'b00110111;
   // assign rom_data[19989]=8'b01010111;
   // assign rom_data[19990]=8'b00110111;
   // assign rom_data[19991]=8'b01010101;
   // assign rom_data[19992]=8'b00110111;
   // assign rom_data[19993]=8'b01010100;
   // assign rom_data[19994]=8'b00110111;
   // assign rom_data[19995]=8'b01010010;
   // assign rom_data[19996]=8'b00110111;
   // assign rom_data[19997]=8'b01010001;
   // assign rom_data[19998]=8'b00110111;
   // assign rom_data[19999]=8'b01010000;
   // assign rom_data[20000]=8'b00110111;
   // assign rom_data[20001]=8'b01001110;
   // assign rom_data[20002]=8'b00110111;
   // assign rom_data[20003]=8'b01001101;
   // assign rom_data[20004]=8'b00110111;
   // assign rom_data[20005]=8'b01001100;
   // assign rom_data[20006]=8'b00110111;
   // assign rom_data[20007]=8'b01001010;
   // assign rom_data[20008]=8'b00110111;
   // assign rom_data[20009]=8'b01001001;
   // assign rom_data[20010]=8'b00110111;
   // assign rom_data[20011]=8'b01000111;
   // assign rom_data[20012]=8'b00110111;
   // assign rom_data[20013]=8'b01000110;
   // assign rom_data[20014]=8'b00110111;
   // assign rom_data[20015]=8'b01000101;
   // assign rom_data[20016]=8'b00110111;
   // assign rom_data[20017]=8'b01000100;
   // assign rom_data[20018]=8'b00110111;
   // assign rom_data[20019]=8'b01000010;
   // assign rom_data[20020]=8'b00110111;
   // assign rom_data[20021]=8'b01000001;
   // assign rom_data[20022]=8'b00110111;
   // assign rom_data[20023]=8'b01000000;
   // assign rom_data[20024]=8'b00110111;
   // assign rom_data[20025]=8'b00111110;
   // assign rom_data[20026]=8'b00110111;
   // assign rom_data[20027]=8'b00111101;
   // assign rom_data[20028]=8'b00110111;
   // assign rom_data[20029]=8'b00111100;
   // assign rom_data[20030]=8'b00110111;
   // assign rom_data[20031]=8'b00111011;
   // assign rom_data[20032]=8'b00110111;
   // assign rom_data[20033]=8'b00111010;
   // assign rom_data[20034]=8'b00110111;
   // assign rom_data[20035]=8'b00111001;
   // assign rom_data[20036]=8'b00110111;
   // assign rom_data[20037]=8'b00110111;
   // assign rom_data[20038]=8'b00110111;
   // assign rom_data[20039]=8'b00110110;
   // assign rom_data[20040]=8'b00110111;
   // assign rom_data[20041]=8'b00110101;
   // assign rom_data[20042]=8'b00110111;
   // assign rom_data[20043]=8'b00110100;
   // assign rom_data[20044]=8'b00110111;
   // assign rom_data[20045]=8'b00110011;
   // assign rom_data[20046]=8'b00110111;
   // assign rom_data[20047]=8'b00110010;
   // assign rom_data[20048]=8'b00110111;
   // assign rom_data[20049]=8'b00110010;
   // assign rom_data[20050]=8'b00110111;
   // assign rom_data[20051]=8'b00110001;
   // assign rom_data[20052]=8'b00110111;
   // assign rom_data[20053]=8'b00110000;
   // assign rom_data[20054]=8'b00110111;
   // assign rom_data[20055]=8'b00101111;
   // assign rom_data[20056]=8'b00110111;
   // assign rom_data[20057]=8'b00101111;
   // assign rom_data[20058]=8'b00110110;
   // assign rom_data[20059]=8'b00101110;
   // assign rom_data[20060]=8'b00110110;
   // assign rom_data[20061]=8'b00101110;
   // assign rom_data[20062]=8'b00110110;
   // assign rom_data[20063]=8'b00101101;
   // assign rom_data[20064]=8'b00110110;
   // assign rom_data[20065]=8'b00101101;
   // assign rom_data[20066]=8'b00110110;
   // assign rom_data[20067]=8'b00101100;
   // assign rom_data[20068]=8'b00110110;
   // assign rom_data[20069]=8'b00101100;
   // assign rom_data[20070]=8'b00110110;
   // assign rom_data[20071]=8'b00101100;
   // assign rom_data[20072]=8'b00110110;
   // assign rom_data[20073]=8'b00101100;
   // assign rom_data[20074]=8'b00110110;
   // assign rom_data[20075]=8'b00101100;
   // assign rom_data[20076]=8'b00110110;
   // assign rom_data[20077]=8'b00101100;
   // assign rom_data[20078]=8'b00110110;
   // assign rom_data[20079]=8'b00101100;
   // assign rom_data[20080]=8'b00110110;
   // assign rom_data[20081]=8'b00101101;
   // assign rom_data[20082]=8'b00110110;
   // assign rom_data[20083]=8'b00101101;
   // assign rom_data[20084]=8'b00110110;
   // assign rom_data[20085]=8'b00101101;
   // assign rom_data[20086]=8'b00110110;
   // assign rom_data[20087]=8'b00101110;
   // assign rom_data[20088]=8'b00110110;
   // assign rom_data[20089]=8'b00101111;
   // assign rom_data[20090]=8'b00110110;
   // assign rom_data[20091]=8'b00101111;
   // assign rom_data[20092]=8'b00110110;
   // assign rom_data[20093]=8'b00110000;
   // assign rom_data[20094]=8'b00110110;
   // assign rom_data[20095]=8'b00110001;
   // assign rom_data[20096]=8'b00110110;
   // assign rom_data[20097]=8'b00110010;
   // assign rom_data[20098]=8'b00110110;
   // assign rom_data[20099]=8'b00110010;
   // assign rom_data[20100]=8'b00110110;
   // assign rom_data[20101]=8'b00110011;
   // assign rom_data[20102]=8'b00110110;
   // assign rom_data[20103]=8'b00110100;
   // assign rom_data[20104]=8'b00110110;
   // assign rom_data[20105]=8'b00110101;
   // assign rom_data[20106]=8'b00110110;
   // assign rom_data[20107]=8'b00110110;
   // assign rom_data[20108]=8'b00110110;
   // assign rom_data[20109]=8'b00110111;
   // assign rom_data[20110]=8'b00110110;
   // assign rom_data[20111]=8'b00111001;
   // assign rom_data[20112]=8'b00110110;
   // assign rom_data[20113]=8'b00111010;
   // assign rom_data[20114]=8'b00110110;
   // assign rom_data[20115]=8'b00111011;
   // assign rom_data[20116]=8'b00110110;
   // assign rom_data[20117]=8'b00111100;
   // assign rom_data[20118]=8'b00110110;
   // assign rom_data[20119]=8'b00111101;
   // assign rom_data[20120]=8'b00110110;
   // assign rom_data[20121]=8'b00111110;
   // assign rom_data[20122]=8'b00110110;
   // assign rom_data[20123]=8'b01000000;
   // assign rom_data[20124]=8'b00110110;
   // assign rom_data[20125]=8'b01000001;
   // assign rom_data[20126]=8'b00110110;
   // assign rom_data[20127]=8'b01000010;
   // assign rom_data[20128]=8'b00110110;
   // assign rom_data[20129]=8'b01000100;
   // assign rom_data[20130]=8'b00110110;
   // assign rom_data[20131]=8'b01000101;
   // assign rom_data[20132]=8'b00110110;
   // assign rom_data[20133]=8'b01000110;
   // assign rom_data[20134]=8'b00110110;
   // assign rom_data[20135]=8'b01001000;
   // assign rom_data[20136]=8'b00110110;
   // assign rom_data[20137]=8'b01001001;
   // assign rom_data[20138]=8'b00110110;
   // assign rom_data[20139]=8'b01001010;
   // assign rom_data[20140]=8'b00110110;
   // assign rom_data[20141]=8'b01001100;
   // assign rom_data[20142]=8'b00110110;
   // assign rom_data[20143]=8'b01001101;
   // assign rom_data[20144]=8'b00110110;
   // assign rom_data[20145]=8'b01001110;
   // assign rom_data[20146]=8'b00110110;
   // assign rom_data[20147]=8'b01010000;
   // assign rom_data[20148]=8'b00110110;
   // assign rom_data[20149]=8'b01010001;
   // assign rom_data[20150]=8'b00110110;
   // assign rom_data[20151]=8'b01010011;
   // assign rom_data[20152]=8'b00110110;
   // assign rom_data[20153]=8'b01010100;
   // assign rom_data[20154]=8'b00110110;
   // assign rom_data[20155]=8'b01010101;
   // assign rom_data[20156]=8'b00110110;
   // assign rom_data[20157]=8'b01010111;
   // assign rom_data[20158]=8'b00110110;
   // assign rom_data[20159]=8'b01011000;
   // assign rom_data[20160]=8'b00110110;
   // assign rom_data[20161]=8'b01011010;
   // assign rom_data[20162]=8'b00110110;
   // assign rom_data[20163]=8'b01011011;
   // assign rom_data[20164]=8'b00110110;
   // assign rom_data[20165]=8'b01011100;
   // assign rom_data[20166]=8'b00110110;
   // assign rom_data[20167]=8'b01011110;
   // assign rom_data[20168]=8'b00110110;
   // assign rom_data[20169]=8'b01011111;
   // assign rom_data[20170]=8'b00110101;
   // assign rom_data[20171]=8'b01100001;
   // assign rom_data[20172]=8'b00110101;
   // assign rom_data[20173]=8'b01100010;
   // assign rom_data[20174]=8'b00110101;
   // assign rom_data[20175]=8'b01100011;
   // assign rom_data[20176]=8'b00110101;
   // assign rom_data[20177]=8'b01100101;
   // assign rom_data[20178]=8'b00110101;
   // assign rom_data[20179]=8'b01100110;
   // assign rom_data[20180]=8'b00110101;
   // assign rom_data[20181]=8'b01101000;
   // assign rom_data[20182]=8'b00110101;
   // assign rom_data[20183]=8'b01101001;
   // assign rom_data[20184]=8'b00110101;
   // assign rom_data[20185]=8'b01101010;
   // assign rom_data[20186]=8'b00110101;
   // assign rom_data[20187]=8'b01101100;
   // assign rom_data[20188]=8'b00110101;
   // assign rom_data[20189]=8'b01101101;
   // assign rom_data[20190]=8'b00110101;
   // assign rom_data[20191]=8'b01101110;
   // assign rom_data[20192]=8'b00110101;
   // assign rom_data[20193]=8'b01110000;
   // assign rom_data[20194]=8'b00110101;
   // assign rom_data[20195]=8'b01110001;
   // assign rom_data[20196]=8'b00110101;
   // assign rom_data[20197]=8'b01110010;
   // assign rom_data[20198]=8'b00110101;
   // assign rom_data[20199]=8'b01110100;
   // assign rom_data[20200]=8'b00110101;
   // assign rom_data[20201]=8'b01110101;
   // assign rom_data[20202]=8'b00110101;
   // assign rom_data[20203]=8'b01110110;
   // assign rom_data[20204]=8'b00110101;
   // assign rom_data[20205]=8'b01110111;
   // assign rom_data[20206]=8'b00110101;
   // assign rom_data[20207]=8'b01111001;
   // assign rom_data[20208]=8'b00110101;
   // assign rom_data[20209]=8'b01111010;
   // assign rom_data[20210]=8'b00110101;
   // assign rom_data[20211]=8'b01111011;
   // assign rom_data[20212]=8'b00110101;
   // assign rom_data[20213]=8'b01111100;
   // assign rom_data[20214]=8'b00110101;
   // assign rom_data[20215]=8'b01111101;
   // assign rom_data[20216]=8'b00110101;
   // assign rom_data[20217]=8'b01111110;
   // assign rom_data[20218]=8'b00110101;
   // assign rom_data[20219]=8'b01111111;
   // assign rom_data[20220]=8'b00110101;
   // assign rom_data[20221]=8'b10000000;
   // assign rom_data[20222]=8'b00110101;
   // assign rom_data[20223]=8'b10000001;
   // assign rom_data[20224]=8'b00110101;
   // assign rom_data[20225]=8'b10000010;
   // assign rom_data[20226]=8'b00110101;
   // assign rom_data[20227]=8'b10000011;
   // assign rom_data[20228]=8'b00110101;
   // assign rom_data[20229]=8'b10000100;
   // assign rom_data[20230]=8'b00110101;
   // assign rom_data[20231]=8'b10000101;
   // assign rom_data[20232]=8'b00110101;
   // assign rom_data[20233]=8'b10000110;
   // assign rom_data[20234]=8'b00110101;
   // assign rom_data[20235]=8'b10000110;
   // assign rom_data[20236]=8'b00110101;
   // assign rom_data[20237]=8'b10000111;
   // assign rom_data[20238]=8'b00110101;
   // assign rom_data[20239]=8'b10001000;
   // assign rom_data[20240]=8'b00110101;
   // assign rom_data[20241]=8'b10001000;
   // assign rom_data[20242]=8'b00110101;
   // assign rom_data[20243]=8'b10001001;
   // assign rom_data[20244]=8'b00110101;
   // assign rom_data[20245]=8'b10001001;
   // assign rom_data[20246]=8'b00110101;
   // assign rom_data[20247]=8'b10001001;
   // assign rom_data[20248]=8'b00110101;
   // assign rom_data[20249]=8'b10001010;
   // assign rom_data[20250]=8'b00110101;
   // assign rom_data[20251]=8'b10001010;
   // assign rom_data[20252]=8'b00110101;
   // assign rom_data[20253]=8'b10001010;
   // assign rom_data[20254]=8'b00110101;
   // assign rom_data[20255]=8'b10001010;
   // assign rom_data[20256]=8'b00110101;
   // assign rom_data[20257]=8'b10001010;
   // assign rom_data[20258]=8'b00110101;
   // assign rom_data[20259]=8'b10001001;
   // assign rom_data[20260]=8'b00110101;
   // assign rom_data[20261]=8'b10001001;
   // assign rom_data[20262]=8'b00110101;
   // assign rom_data[20263]=8'b10001001;
   // assign rom_data[20264]=8'b00110101;
   // assign rom_data[20265]=8'b10001000;
   // assign rom_data[20266]=8'b00110101;
   // assign rom_data[20267]=8'b10001000;
   // assign rom_data[20268]=8'b00110101;
   // assign rom_data[20269]=8'b10000111;
   // assign rom_data[20270]=8'b00110101;
   // assign rom_data[20271]=8'b10000111;
   // assign rom_data[20272]=8'b00110101;
   // assign rom_data[20273]=8'b10000110;
   // assign rom_data[20274]=8'b00110101;
   // assign rom_data[20275]=8'b10000101;
   // assign rom_data[20276]=8'b00110101;
   // assign rom_data[20277]=8'b10000100;
   // assign rom_data[20278]=8'b00110100;
   // assign rom_data[20279]=8'b10000011;
   // assign rom_data[20280]=8'b00110100;
   // assign rom_data[20281]=8'b10000010;
   // assign rom_data[20282]=8'b00110100;
   // assign rom_data[20283]=8'b10000010;
   // assign rom_data[20284]=8'b00110100;
   // assign rom_data[20285]=8'b10000001;
   // assign rom_data[20286]=8'b00110100;
   // assign rom_data[20287]=8'b01111111;
   // assign rom_data[20288]=8'b00110100;
   // assign rom_data[20289]=8'b01111110;
   // assign rom_data[20290]=8'b00110100;
   // assign rom_data[20291]=8'b01111101;
   // assign rom_data[20292]=8'b00110100;
   // assign rom_data[20293]=8'b01111100;
   // assign rom_data[20294]=8'b00110100;
   // assign rom_data[20295]=8'b01111011;
   // assign rom_data[20296]=8'b00110100;
   // assign rom_data[20297]=8'b01111010;
   // assign rom_data[20298]=8'b00110100;
   // assign rom_data[20299]=8'b01111001;
   // assign rom_data[20300]=8'b00110100;
   // assign rom_data[20301]=8'b01110111;
   // assign rom_data[20302]=8'b00110100;
   // assign rom_data[20303]=8'b01110110;
   // assign rom_data[20304]=8'b00110100;
   // assign rom_data[20305]=8'b01110101;
   // assign rom_data[20306]=8'b00110100;
   // assign rom_data[20307]=8'b01110100;
   // assign rom_data[20308]=8'b00110100;
   // assign rom_data[20309]=8'b01110010;
   // assign rom_data[20310]=8'b00110100;
   // assign rom_data[20311]=8'b01110001;
   // assign rom_data[20312]=8'b00110100;
   // assign rom_data[20313]=8'b01110000;
   // assign rom_data[20314]=8'b00110100;
   // assign rom_data[20315]=8'b01101110;
   // assign rom_data[20316]=8'b00110100;
   // assign rom_data[20317]=8'b01101101;
   // assign rom_data[20318]=8'b00110100;
   // assign rom_data[20319]=8'b01101100;
   // assign rom_data[20320]=8'b00110100;
   // assign rom_data[20321]=8'b01101010;
   // assign rom_data[20322]=8'b00110100;
   // assign rom_data[20323]=8'b01101001;
   // assign rom_data[20324]=8'b00110100;
   // assign rom_data[20325]=8'b01100111;
   // assign rom_data[20326]=8'b00110100;
   // assign rom_data[20327]=8'b01100110;
   // assign rom_data[20328]=8'b00110100;
   // assign rom_data[20329]=8'b01100101;
   // assign rom_data[20330]=8'b00110100;
   // assign rom_data[20331]=8'b01100011;
   // assign rom_data[20332]=8'b00110100;
   // assign rom_data[20333]=8'b01100010;
   // assign rom_data[20334]=8'b00110100;
   // assign rom_data[20335]=8'b01100000;
   // assign rom_data[20336]=8'b00110100;
   // assign rom_data[20337]=8'b01011111;
   // assign rom_data[20338]=8'b00110100;
   // assign rom_data[20339]=8'b01011110;
   // assign rom_data[20340]=8'b00110100;
   // assign rom_data[20341]=8'b01011100;
   // assign rom_data[20342]=8'b00110100;
   // assign rom_data[20343]=8'b01011011;
   // assign rom_data[20344]=8'b00110100;
   // assign rom_data[20345]=8'b01011001;
   // assign rom_data[20346]=8'b00110100;
   // assign rom_data[20347]=8'b01011000;
   // assign rom_data[20348]=8'b00110100;
   // assign rom_data[20349]=8'b01010111;
   // assign rom_data[20350]=8'b00110100;
   // assign rom_data[20351]=8'b01010101;
   // assign rom_data[20352]=8'b00110100;
   // assign rom_data[20353]=8'b01010100;
   // assign rom_data[20354]=8'b00110100;
   // assign rom_data[20355]=8'b01010010;
   // assign rom_data[20356]=8'b00110100;
   // assign rom_data[20357]=8'b01010001;
   // assign rom_data[20358]=8'b00110100;
   // assign rom_data[20359]=8'b01010000;
   // assign rom_data[20360]=8'b00110100;
   // assign rom_data[20361]=8'b01001110;
   // assign rom_data[20362]=8'b00110100;
   // assign rom_data[20363]=8'b01001101;
   // assign rom_data[20364]=8'b00110100;
   // assign rom_data[20365]=8'b01001011;
   // assign rom_data[20366]=8'b00110100;
   // assign rom_data[20367]=8'b01001010;
   // assign rom_data[20368]=8'b00110100;
   // assign rom_data[20369]=8'b01001001;
   // assign rom_data[20370]=8'b00110100;
   // assign rom_data[20371]=8'b01000111;
   // assign rom_data[20372]=8'b00110100;
   // assign rom_data[20373]=8'b01000110;
   // assign rom_data[20374]=8'b00110100;
   // assign rom_data[20375]=8'b01000101;
   // assign rom_data[20376]=8'b00110100;
   // assign rom_data[20377]=8'b01000011;
   // assign rom_data[20378]=8'b00110100;
   // assign rom_data[20379]=8'b01000010;
   // assign rom_data[20380]=8'b00110100;
   // assign rom_data[20381]=8'b01000001;
   // assign rom_data[20382]=8'b00110100;
   // assign rom_data[20383]=8'b01000000;
   // assign rom_data[20384]=8'b00110100;
   // assign rom_data[20385]=8'b00111110;
   // assign rom_data[20386]=8'b00110100;
   // assign rom_data[20387]=8'b00111101;
   // assign rom_data[20388]=8'b00110100;
   // assign rom_data[20389]=8'b00111100;
   // assign rom_data[20390]=8'b00110100;
   // assign rom_data[20391]=8'b00111011;
   // assign rom_data[20392]=8'b00110100;
   // assign rom_data[20393]=8'b00111010;
   // assign rom_data[20394]=8'b00110100;
   // assign rom_data[20395]=8'b00111001;
   // assign rom_data[20396]=8'b00110100;
   // assign rom_data[20397]=8'b00110111;
   // assign rom_data[20398]=8'b00110100;
   // assign rom_data[20399]=8'b00110110;
   // assign rom_data[20400]=8'b00110011;
   // assign rom_data[20401]=8'b00110101;
   // assign rom_data[20402]=8'b00110011;
   // assign rom_data[20403]=8'b00110100;
   // assign rom_data[20404]=8'b00110011;
   // assign rom_data[20405]=8'b00110011;
   // assign rom_data[20406]=8'b00110011;
   // assign rom_data[20407]=8'b00110010;
   // assign rom_data[20408]=8'b00110011;
   // assign rom_data[20409]=8'b00110010;
   // assign rom_data[20410]=8'b00110011;
   // assign rom_data[20411]=8'b00110001;
   // assign rom_data[20412]=8'b00110011;
   // assign rom_data[20413]=8'b00110000;
   // assign rom_data[20414]=8'b00110011;
   // assign rom_data[20415]=8'b00101111;
   // assign rom_data[20416]=8'b00110011;
   // assign rom_data[20417]=8'b00101111;
   // assign rom_data[20418]=8'b00110011;
   // assign rom_data[20419]=8'b00101110;
   // assign rom_data[20420]=8'b00110011;
   // assign rom_data[20421]=8'b00101110;
   // assign rom_data[20422]=8'b00110011;
   // assign rom_data[20423]=8'b00101101;
   // assign rom_data[20424]=8'b00110011;
   // assign rom_data[20425]=8'b00101101;
   // assign rom_data[20426]=8'b00110011;
   // assign rom_data[20427]=8'b00101100;
   // assign rom_data[20428]=8'b00110011;
   // assign rom_data[20429]=8'b00101100;
   // assign rom_data[20430]=8'b00110011;
   // assign rom_data[20431]=8'b00101100;
   // assign rom_data[20432]=8'b00110011;
   // assign rom_data[20433]=8'b00101100;
   // assign rom_data[20434]=8'b00110011;
   // assign rom_data[20435]=8'b00101100;
   // assign rom_data[20436]=8'b00110011;
   // assign rom_data[20437]=8'b00101100;
   // assign rom_data[20438]=8'b00110011;
   // assign rom_data[20439]=8'b00101100;
   // assign rom_data[20440]=8'b00110011;
   // assign rom_data[20441]=8'b00101101;
   // assign rom_data[20442]=8'b00110011;
   // assign rom_data[20443]=8'b00101101;
   // assign rom_data[20444]=8'b00110011;
   // assign rom_data[20445]=8'b00101101;
   // assign rom_data[20446]=8'b00110011;
   // assign rom_data[20447]=8'b00101110;
   // assign rom_data[20448]=8'b00110011;
   // assign rom_data[20449]=8'b00101111;
   // assign rom_data[20450]=8'b00110011;
   // assign rom_data[20451]=8'b00101111;
   // assign rom_data[20452]=8'b00110011;
   // assign rom_data[20453]=8'b00110000;
   // assign rom_data[20454]=8'b00110011;
   // assign rom_data[20455]=8'b00110001;
   // assign rom_data[20456]=8'b00110011;
   // assign rom_data[20457]=8'b00110010;
   // assign rom_data[20458]=8'b00110011;
   // assign rom_data[20459]=8'b00110010;
   // assign rom_data[20460]=8'b00110011;
   // assign rom_data[20461]=8'b00110011;
   // assign rom_data[20462]=8'b00110011;
   // assign rom_data[20463]=8'b00110100;
   // assign rom_data[20464]=8'b00110011;
   // assign rom_data[20465]=8'b00110101;
   // assign rom_data[20466]=8'b00110011;
   // assign rom_data[20467]=8'b00110110;
   // assign rom_data[20468]=8'b00110011;
   // assign rom_data[20469]=8'b00110111;
   // assign rom_data[20470]=8'b00110011;
   // assign rom_data[20471]=8'b00111001;
   // assign rom_data[20472]=8'b00110011;
   // assign rom_data[20473]=8'b00111010;
   // assign rom_data[20474]=8'b00110011;
   // assign rom_data[20475]=8'b00111011;
   // assign rom_data[20476]=8'b00110011;
   // assign rom_data[20477]=8'b00111100;
   // assign rom_data[20478]=8'b00110011;
   // assign rom_data[20479]=8'b00111101;
   // assign rom_data[20480]=8'b00110011;
   // assign rom_data[20481]=8'b00111110;
   // assign rom_data[20482]=8'b00110011;
   // assign rom_data[20483]=8'b01000000;
   // assign rom_data[20484]=8'b00110011;
   // assign rom_data[20485]=8'b01000001;
   // assign rom_data[20486]=8'b00110011;
   // assign rom_data[20487]=8'b01000010;
   // assign rom_data[20488]=8'b00110011;
   // assign rom_data[20489]=8'b01000100;
   // assign rom_data[20490]=8'b00110011;
   // assign rom_data[20491]=8'b01000101;
   // assign rom_data[20492]=8'b00110011;
   // assign rom_data[20493]=8'b01000110;
   // assign rom_data[20494]=8'b00110011;
   // assign rom_data[20495]=8'b01001000;
   // assign rom_data[20496]=8'b00110011;
   // assign rom_data[20497]=8'b01001001;
   // assign rom_data[20498]=8'b00110011;
   // assign rom_data[20499]=8'b01001010;
   // assign rom_data[20500]=8'b00110011;
   // assign rom_data[20501]=8'b01001100;
   // assign rom_data[20502]=8'b00110011;
   // assign rom_data[20503]=8'b01001101;
   // assign rom_data[20504]=8'b00110011;
   // assign rom_data[20505]=8'b01001110;
   // assign rom_data[20506]=8'b00110010;
   // assign rom_data[20507]=8'b01010000;
   // assign rom_data[20508]=8'b00110010;
   // assign rom_data[20509]=8'b01010001;
   // assign rom_data[20510]=8'b00110010;
   // assign rom_data[20511]=8'b01010011;
   // assign rom_data[20512]=8'b00110010;
   // assign rom_data[20513]=8'b01010100;
   // assign rom_data[20514]=8'b00110010;
   // assign rom_data[20515]=8'b01010101;
   // assign rom_data[20516]=8'b00110010;
   // assign rom_data[20517]=8'b01010111;
   // assign rom_data[20518]=8'b00110010;
   // assign rom_data[20519]=8'b01011000;
   // assign rom_data[20520]=8'b00110010;
   // assign rom_data[20521]=8'b01011010;
   // assign rom_data[20522]=8'b00110010;
   // assign rom_data[20523]=8'b01011011;
   // assign rom_data[20524]=8'b00110010;
   // assign rom_data[20525]=8'b01011100;
   // assign rom_data[20526]=8'b00110010;
   // assign rom_data[20527]=8'b01011110;
   // assign rom_data[20528]=8'b00110010;
   // assign rom_data[20529]=8'b01011111;
   // assign rom_data[20530]=8'b00110010;
   // assign rom_data[20531]=8'b01100001;
   // assign rom_data[20532]=8'b00110010;
   // assign rom_data[20533]=8'b01100010;
   // assign rom_data[20534]=8'b00110010;
   // assign rom_data[20535]=8'b01100011;
   // assign rom_data[20536]=8'b00110010;
   // assign rom_data[20537]=8'b01100101;
   // assign rom_data[20538]=8'b00110010;
   // assign rom_data[20539]=8'b01100110;
   // assign rom_data[20540]=8'b00110010;
   // assign rom_data[20541]=8'b01101000;
   // assign rom_data[20542]=8'b00110010;
   // assign rom_data[20543]=8'b01101001;
   // assign rom_data[20544]=8'b00110010;
   // assign rom_data[20545]=8'b01101010;
   // assign rom_data[20546]=8'b00110010;
   // assign rom_data[20547]=8'b01101100;
   // assign rom_data[20548]=8'b00110010;
   // assign rom_data[20549]=8'b01101101;
   // assign rom_data[20550]=8'b00110010;
   // assign rom_data[20551]=8'b01101110;
   // assign rom_data[20552]=8'b00110010;
   // assign rom_data[20553]=8'b01110000;
   // assign rom_data[20554]=8'b00110010;
   // assign rom_data[20555]=8'b01110001;
   // assign rom_data[20556]=8'b00110010;
   // assign rom_data[20557]=8'b01110010;
   // assign rom_data[20558]=8'b00110010;
   // assign rom_data[20559]=8'b01110100;
   // assign rom_data[20560]=8'b00110010;
   // assign rom_data[20561]=8'b01110101;
   // assign rom_data[20562]=8'b00110010;
   // assign rom_data[20563]=8'b01110110;
   // assign rom_data[20564]=8'b00110010;
   // assign rom_data[20565]=8'b01110111;
   // assign rom_data[20566]=8'b00110010;
   // assign rom_data[20567]=8'b01111001;
   // assign rom_data[20568]=8'b00110010;
   // assign rom_data[20569]=8'b01111010;
   // assign rom_data[20570]=8'b00110010;
   // assign rom_data[20571]=8'b01111011;
   // assign rom_data[20572]=8'b00110010;
   // assign rom_data[20573]=8'b01111100;
   // assign rom_data[20574]=8'b00110010;
   // assign rom_data[20575]=8'b01111101;
   // assign rom_data[20576]=8'b00110010;
   // assign rom_data[20577]=8'b01111110;
   // assign rom_data[20578]=8'b00110010;
   // assign rom_data[20579]=8'b01111111;
   // assign rom_data[20580]=8'b00110010;
   // assign rom_data[20581]=8'b10000000;
   // assign rom_data[20582]=8'b00110010;
   // assign rom_data[20583]=8'b10000001;
   // assign rom_data[20584]=8'b00110010;
   // assign rom_data[20585]=8'b10000010;
   // assign rom_data[20586]=8'b00110010;
   // assign rom_data[20587]=8'b10000011;
   // assign rom_data[20588]=8'b00110010;
   // assign rom_data[20589]=8'b10000100;
   // assign rom_data[20590]=8'b00110010;
   // assign rom_data[20591]=8'b10000101;
   // assign rom_data[20592]=8'b00110010;
   // assign rom_data[20593]=8'b10000110;
   // assign rom_data[20594]=8'b00110010;
   // assign rom_data[20595]=8'b10000111;
   // assign rom_data[20596]=8'b00110010;
   // assign rom_data[20597]=8'b10000111;
   // assign rom_data[20598]=8'b00110010;
   // assign rom_data[20599]=8'b10001000;
   // assign rom_data[20600]=8'b00110010;
   // assign rom_data[20601]=8'b10001000;
   // assign rom_data[20602]=8'b00110010;
   // assign rom_data[20603]=8'b10001001;
   // assign rom_data[20604]=8'b00110010;
   // assign rom_data[20605]=8'b10001001;
   // assign rom_data[20606]=8'b00110010;
   // assign rom_data[20607]=8'b10001001;
   // assign rom_data[20608]=8'b00110010;
   // assign rom_data[20609]=8'b10001010;
   // assign rom_data[20610]=8'b00110010;
   // assign rom_data[20611]=8'b10001010;
   // assign rom_data[20612]=8'b00110010;
   // assign rom_data[20613]=8'b10001010;
   // assign rom_data[20614]=8'b00110010;
   // assign rom_data[20615]=8'b10001010;
   // assign rom_data[20616]=8'b00110010;
   // assign rom_data[20617]=8'b10001010;
   // assign rom_data[20618]=8'b00110010;
   // assign rom_data[20619]=8'b10001001;
   // assign rom_data[20620]=8'b00110001;
   // assign rom_data[20621]=8'b10001001;
   // assign rom_data[20622]=8'b00110001;
   // assign rom_data[20623]=8'b10001001;
   // assign rom_data[20624]=8'b00110001;
   // assign rom_data[20625]=8'b10001000;
   // assign rom_data[20626]=8'b00110001;
   // assign rom_data[20627]=8'b10001000;
   // assign rom_data[20628]=8'b00110001;
   // assign rom_data[20629]=8'b10000111;
   // assign rom_data[20630]=8'b00110001;
   // assign rom_data[20631]=8'b10000111;
   // assign rom_data[20632]=8'b00110001;
   // assign rom_data[20633]=8'b10000110;
   // assign rom_data[20634]=8'b00110001;
   // assign rom_data[20635]=8'b10000101;
   // assign rom_data[20636]=8'b00110001;
   // assign rom_data[20637]=8'b10000100;
   // assign rom_data[20638]=8'b00110001;
   // assign rom_data[20639]=8'b10000011;
   // assign rom_data[20640]=8'b00110001;
   // assign rom_data[20641]=8'b10000010;
   // assign rom_data[20642]=8'b00110001;
   // assign rom_data[20643]=8'b10000010;
   // assign rom_data[20644]=8'b00110001;
   // assign rom_data[20645]=8'b10000001;
   // assign rom_data[20646]=8'b00110001;
   // assign rom_data[20647]=8'b01111111;
   // assign rom_data[20648]=8'b00110001;
   // assign rom_data[20649]=8'b01111110;
   // assign rom_data[20650]=8'b00110001;
   // assign rom_data[20651]=8'b01111101;
   // assign rom_data[20652]=8'b00110001;
   // assign rom_data[20653]=8'b01111100;
   // assign rom_data[20654]=8'b00110001;
   // assign rom_data[20655]=8'b01111011;
   // assign rom_data[20656]=8'b00110001;
   // assign rom_data[20657]=8'b01111010;
   // assign rom_data[20658]=8'b00110001;
   // assign rom_data[20659]=8'b01111001;
   // assign rom_data[20660]=8'b00110001;
   // assign rom_data[20661]=8'b01110111;
   // assign rom_data[20662]=8'b00110001;
   // assign rom_data[20663]=8'b01110110;
   // assign rom_data[20664]=8'b00110001;
   // assign rom_data[20665]=8'b01110101;
   // assign rom_data[20666]=8'b00110001;
   // assign rom_data[20667]=8'b01110100;
   // assign rom_data[20668]=8'b00110001;
   // assign rom_data[20669]=8'b01110010;
   // assign rom_data[20670]=8'b00110001;
   // assign rom_data[20671]=8'b01110001;
   // assign rom_data[20672]=8'b00110001;
   // assign rom_data[20673]=8'b01110000;
   // assign rom_data[20674]=8'b00110001;
   // assign rom_data[20675]=8'b01101110;
   // assign rom_data[20676]=8'b00110001;
   // assign rom_data[20677]=8'b01101101;
   // assign rom_data[20678]=8'b00110001;
   // assign rom_data[20679]=8'b01101100;
   // assign rom_data[20680]=8'b00110001;
   // assign rom_data[20681]=8'b01101010;
   // assign rom_data[20682]=8'b00110001;
   // assign rom_data[20683]=8'b01101001;
   // assign rom_data[20684]=8'b00110001;
   // assign rom_data[20685]=8'b01100111;
   // assign rom_data[20686]=8'b00110001;
   // assign rom_data[20687]=8'b01100110;
   // assign rom_data[20688]=8'b00110001;
   // assign rom_data[20689]=8'b01100101;
   // assign rom_data[20690]=8'b00110001;
   // assign rom_data[20691]=8'b01100011;
   // assign rom_data[20692]=8'b00110001;
   // assign rom_data[20693]=8'b01100010;
   // assign rom_data[20694]=8'b00110001;
   // assign rom_data[20695]=8'b01100000;
   // assign rom_data[20696]=8'b00110001;
   // assign rom_data[20697]=8'b01011111;
   // assign rom_data[20698]=8'b00110001;
   // assign rom_data[20699]=8'b01011110;
   // assign rom_data[20700]=8'b00110001;
   // assign rom_data[20701]=8'b01011100;
   // assign rom_data[20702]=8'b00110001;
   // assign rom_data[20703]=8'b01011011;
   // assign rom_data[20704]=8'b00110001;
   // assign rom_data[20705]=8'b01011001;
   // assign rom_data[20706]=8'b00110001;
   // assign rom_data[20707]=8'b01011000;
   // assign rom_data[20708]=8'b00110001;
   // assign rom_data[20709]=8'b01010111;
   // assign rom_data[20710]=8'b00110001;
   // assign rom_data[20711]=8'b01010101;
   // assign rom_data[20712]=8'b00110001;
   // assign rom_data[20713]=8'b01010100;
   // assign rom_data[20714]=8'b00110001;
   // assign rom_data[20715]=8'b01010010;
   // assign rom_data[20716]=8'b00110001;
   // assign rom_data[20717]=8'b01010001;
   // assign rom_data[20718]=8'b00110001;
   // assign rom_data[20719]=8'b01010000;
   // assign rom_data[20720]=8'b00110001;
   // assign rom_data[20721]=8'b01001110;
   // assign rom_data[20722]=8'b00110001;
   // assign rom_data[20723]=8'b01001101;
   // assign rom_data[20724]=8'b00110001;
   // assign rom_data[20725]=8'b01001011;
   // assign rom_data[20726]=8'b00110001;
   // assign rom_data[20727]=8'b01001010;
   // assign rom_data[20728]=8'b00110001;
   // assign rom_data[20729]=8'b01001001;
   // assign rom_data[20730]=8'b00110001;
   // assign rom_data[20731]=8'b01000111;
   // assign rom_data[20732]=8'b00110001;
   // assign rom_data[20733]=8'b01000110;
   // assign rom_data[20734]=8'b00110001;
   // assign rom_data[20735]=8'b01000101;
   // assign rom_data[20736]=8'b00110001;
   // assign rom_data[20737]=8'b01000011;
   // assign rom_data[20738]=8'b00110001;
   // assign rom_data[20739]=8'b01000010;
   // assign rom_data[20740]=8'b00110000;
   // assign rom_data[20741]=8'b01000001;
   // assign rom_data[20742]=8'b00110000;
   // assign rom_data[20743]=8'b01000000;
   // assign rom_data[20744]=8'b00110000;
   // assign rom_data[20745]=8'b00111110;
   // assign rom_data[20746]=8'b00110000;
   // assign rom_data[20747]=8'b00111101;
   // assign rom_data[20748]=8'b00110000;
   // assign rom_data[20749]=8'b00111100;
   // assign rom_data[20750]=8'b00110000;
   // assign rom_data[20751]=8'b00111011;
   // assign rom_data[20752]=8'b00110000;
   // assign rom_data[20753]=8'b00111010;
   // assign rom_data[20754]=8'b00110000;
   // assign rom_data[20755]=8'b00111001;
   // assign rom_data[20756]=8'b00110000;
   // assign rom_data[20757]=8'b00110111;
   // assign rom_data[20758]=8'b00110000;
   // assign rom_data[20759]=8'b00110110;
   // assign rom_data[20760]=8'b00110000;
   // assign rom_data[20761]=8'b00110101;
   // assign rom_data[20762]=8'b00110000;
   // assign rom_data[20763]=8'b00110100;
   // assign rom_data[20764]=8'b00110000;
   // assign rom_data[20765]=8'b00110011;
   // assign rom_data[20766]=8'b00110000;
   // assign rom_data[20767]=8'b00110010;
   // assign rom_data[20768]=8'b00110000;
   // assign rom_data[20769]=8'b00110010;
   // assign rom_data[20770]=8'b00110000;
   // assign rom_data[20771]=8'b00110001;
   // assign rom_data[20772]=8'b00110000;
   // assign rom_data[20773]=8'b00110000;
   // assign rom_data[20774]=8'b00110000;
   // assign rom_data[20775]=8'b00101111;
   // assign rom_data[20776]=8'b00110000;
   // assign rom_data[20777]=8'b00101111;
   // assign rom_data[20778]=8'b00110000;
   // assign rom_data[20779]=8'b00101110;
   // assign rom_data[20780]=8'b00110000;
   // assign rom_data[20781]=8'b00101110;
   // assign rom_data[20782]=8'b00110000;
   // assign rom_data[20783]=8'b00101101;
   // assign rom_data[20784]=8'b00110000;
   // assign rom_data[20785]=8'b00101101;
   // assign rom_data[20786]=8'b00110000;
   // assign rom_data[20787]=8'b00101100;
   // assign rom_data[20788]=8'b00110000;
   // assign rom_data[20789]=8'b00101100;
   // assign rom_data[20790]=8'b00110000;
   // assign rom_data[20791]=8'b00101100;
   // assign rom_data[20792]=8'b00110000;
   // assign rom_data[20793]=8'b00101100;
   // assign rom_data[20794]=8'b00110000;
   // assign rom_data[20795]=8'b00101100;
   // assign rom_data[20796]=8'b00110000;
   // assign rom_data[20797]=8'b00101100;
   // assign rom_data[20798]=8'b00110000;
   // assign rom_data[20799]=8'b00101100;
   // assign rom_data[20800]=8'b00110000;
   // assign rom_data[20801]=8'b00101101;
   // assign rom_data[20802]=8'b00110000;
   // assign rom_data[20803]=8'b00101101;
   // assign rom_data[20804]=8'b00110000;
   // assign rom_data[20805]=8'b00101101;
   // assign rom_data[20806]=8'b00110000;
   // assign rom_data[20807]=8'b00101110;
   // assign rom_data[20808]=8'b00110000;
   // assign rom_data[20809]=8'b00101111;
   // assign rom_data[20810]=8'b00110000;
   // assign rom_data[20811]=8'b00101111;
   // assign rom_data[20812]=8'b00110000;
   // assign rom_data[20813]=8'b00110000;
   // assign rom_data[20814]=8'b00110000;
   // assign rom_data[20815]=8'b00110001;
   // assign rom_data[20816]=8'b00110000;
   // assign rom_data[20817]=8'b00110010;
   // assign rom_data[20818]=8'b00110000;
   // assign rom_data[20819]=8'b00110010;
   // assign rom_data[20820]=8'b00110000;
   // assign rom_data[20821]=8'b00110011;
   // assign rom_data[20822]=8'b00110000;
   // assign rom_data[20823]=8'b00110100;
   // assign rom_data[20824]=8'b00110000;
   // assign rom_data[20825]=8'b00110101;
   // assign rom_data[20826]=8'b00110000;
   // assign rom_data[20827]=8'b00110110;
   // assign rom_data[20828]=8'b00110000;
   // assign rom_data[20829]=8'b00110111;
   // assign rom_data[20830]=8'b00110000;
   // assign rom_data[20831]=8'b00111001;
   // assign rom_data[20832]=8'b00110000;
   // assign rom_data[20833]=8'b00111010;
   // assign rom_data[20834]=8'b00110000;
   // assign rom_data[20835]=8'b00111011;
   // assign rom_data[20836]=8'b00110000;
   // assign rom_data[20837]=8'b00111100;
   // assign rom_data[20838]=8'b00110000;
   // assign rom_data[20839]=8'b00111101;
   // assign rom_data[20840]=8'b00110000;
   // assign rom_data[20841]=8'b00111110;
   // assign rom_data[20842]=8'b00110000;
   // assign rom_data[20843]=8'b01000000;
   // assign rom_data[20844]=8'b00101111;
   // assign rom_data[20845]=8'b01000001;
   // assign rom_data[20846]=8'b00101111;
   // assign rom_data[20847]=8'b01000010;
   // assign rom_data[20848]=8'b00101111;
   // assign rom_data[20849]=8'b01000100;
   // assign rom_data[20850]=8'b00101111;
   // assign rom_data[20851]=8'b01000101;
   // assign rom_data[20852]=8'b00101111;
   // assign rom_data[20853]=8'b01000110;
   // assign rom_data[20854]=8'b00101111;
   // assign rom_data[20855]=8'b01001000;
   // assign rom_data[20856]=8'b00101111;
   // assign rom_data[20857]=8'b01001001;
   // assign rom_data[20858]=8'b00101111;
   // assign rom_data[20859]=8'b01001010;
   // assign rom_data[20860]=8'b00101111;
   // assign rom_data[20861]=8'b01001100;
   // assign rom_data[20862]=8'b00101111;
   // assign rom_data[20863]=8'b01001101;
   // assign rom_data[20864]=8'b00101111;
   // assign rom_data[20865]=8'b01001110;
   // assign rom_data[20866]=8'b00101111;
   // assign rom_data[20867]=8'b01010000;
   // assign rom_data[20868]=8'b00101111;
   // assign rom_data[20869]=8'b01010001;
   // assign rom_data[20870]=8'b00101111;
   // assign rom_data[20871]=8'b01010011;
   // assign rom_data[20872]=8'b00101111;
   // assign rom_data[20873]=8'b01010100;
   // assign rom_data[20874]=8'b00101111;
   // assign rom_data[20875]=8'b01010101;
   // assign rom_data[20876]=8'b00101111;
   // assign rom_data[20877]=8'b01010111;
   // assign rom_data[20878]=8'b00101111;
   // assign rom_data[20879]=8'b01011000;
   // assign rom_data[20880]=8'b00101111;
   // assign rom_data[20881]=8'b01011010;
   // assign rom_data[20882]=8'b00101111;
   // assign rom_data[20883]=8'b01011011;
   // assign rom_data[20884]=8'b00101111;
   // assign rom_data[20885]=8'b01011100;
   // assign rom_data[20886]=8'b00101111;
   // assign rom_data[20887]=8'b01011110;
   // assign rom_data[20888]=8'b00101111;
   // assign rom_data[20889]=8'b01011111;
   // assign rom_data[20890]=8'b00101111;
   // assign rom_data[20891]=8'b01100001;
   // assign rom_data[20892]=8'b00101111;
   // assign rom_data[20893]=8'b01100010;
   // assign rom_data[20894]=8'b00101111;
   // assign rom_data[20895]=8'b01100011;
   // assign rom_data[20896]=8'b00101111;
   // assign rom_data[20897]=8'b01100101;
   // assign rom_data[20898]=8'b00101111;
   // assign rom_data[20899]=8'b01100110;
   // assign rom_data[20900]=8'b00101111;
   // assign rom_data[20901]=8'b01101000;
   // assign rom_data[20902]=8'b00101111;
   // assign rom_data[20903]=8'b01101001;
   // assign rom_data[20904]=8'b00101111;
   // assign rom_data[20905]=8'b01101010;
   // assign rom_data[20906]=8'b00101111;
   // assign rom_data[20907]=8'b01101100;
   // assign rom_data[20908]=8'b00101111;
   // assign rom_data[20909]=8'b01101101;
   // assign rom_data[20910]=8'b00101111;
   // assign rom_data[20911]=8'b01101110;
   // assign rom_data[20912]=8'b00101111;
   // assign rom_data[20913]=8'b01110000;
   // assign rom_data[20914]=8'b00101111;
   // assign rom_data[20915]=8'b01110001;
   // assign rom_data[20916]=8'b00101111;
   // assign rom_data[20917]=8'b01110010;
   // assign rom_data[20918]=8'b00101111;
   // assign rom_data[20919]=8'b01110100;
   // assign rom_data[20920]=8'b00101111;
   // assign rom_data[20921]=8'b01110101;
   // assign rom_data[20922]=8'b00101111;
   // assign rom_data[20923]=8'b01110110;
   // assign rom_data[20924]=8'b00101111;
   // assign rom_data[20925]=8'b01110111;
   // assign rom_data[20926]=8'b00101111;
   // assign rom_data[20927]=8'b01111001;
   // assign rom_data[20928]=8'b00101111;
   // assign rom_data[20929]=8'b01111010;
   // assign rom_data[20930]=8'b00101111;
   // assign rom_data[20931]=8'b01111011;
   // assign rom_data[20932]=8'b00101111;
   // assign rom_data[20933]=8'b01111100;
   // assign rom_data[20934]=8'b00101111;
   // assign rom_data[20935]=8'b01111101;
   // assign rom_data[20936]=8'b00101111;
   // assign rom_data[20937]=8'b01111110;
   // assign rom_data[20938]=8'b00101111;
   // assign rom_data[20939]=8'b01111111;
   // assign rom_data[20940]=8'b00101111;
   // assign rom_data[20941]=8'b10000000;
   // assign rom_data[20942]=8'b00101111;
   // assign rom_data[20943]=8'b10000001;
   // assign rom_data[20944]=8'b00101111;
   // assign rom_data[20945]=8'b10000010;
   // assign rom_data[20946]=8'b00101111;
   // assign rom_data[20947]=8'b10000011;
   // assign rom_data[20948]=8'b00101111;
   // assign rom_data[20949]=8'b10000100;
   // assign rom_data[20950]=8'b00101111;
   // assign rom_data[20951]=8'b10000101;
   // assign rom_data[20952]=8'b00101111;
   // assign rom_data[20953]=8'b10000110;
   // assign rom_data[20954]=8'b00101111;
   // assign rom_data[20955]=8'b10000111;
   // assign rom_data[20956]=8'b00101111;
   // assign rom_data[20957]=8'b10000111;
   // assign rom_data[20958]=8'b00101111;
   // assign rom_data[20959]=8'b10001000;
   // assign rom_data[20960]=8'b00101111;
   // assign rom_data[20961]=8'b10001000;
   // assign rom_data[20962]=8'b00101110;
   // assign rom_data[20963]=8'b10001001;
   // assign rom_data[20964]=8'b00101110;
   // assign rom_data[20965]=8'b10001001;
   // assign rom_data[20966]=8'b00101110;
   // assign rom_data[20967]=8'b10001001;
   // assign rom_data[20968]=8'b00101110;
   // assign rom_data[20969]=8'b10001010;
   // assign rom_data[20970]=8'b00101110;
   // assign rom_data[20971]=8'b10001010;
   // assign rom_data[20972]=8'b00101110;
   // assign rom_data[20973]=8'b10001010;
   // assign rom_data[20974]=8'b00101110;
   // assign rom_data[20975]=8'b10001010;
   // assign rom_data[20976]=8'b00101110;
   // assign rom_data[20977]=8'b10001010;
   // assign rom_data[20978]=8'b00101110;
   // assign rom_data[20979]=8'b10001001;
   // assign rom_data[20980]=8'b00101110;
   // assign rom_data[20981]=8'b10001001;
   // assign rom_data[20982]=8'b00101110;
   // assign rom_data[20983]=8'b10001001;
   // assign rom_data[20984]=8'b00101110;
   // assign rom_data[20985]=8'b10001000;
   // assign rom_data[20986]=8'b00101110;
   // assign rom_data[20987]=8'b10001000;
   // assign rom_data[20988]=8'b00101110;
   // assign rom_data[20989]=8'b10000111;
   // assign rom_data[20990]=8'b00101110;
   // assign rom_data[20991]=8'b10000111;
   // assign rom_data[20992]=8'b00101110;
   // assign rom_data[20993]=8'b10000110;
   // assign rom_data[20994]=8'b00101110;
   // assign rom_data[20995]=8'b10000101;
   // assign rom_data[20996]=8'b00101110;
   // assign rom_data[20997]=8'b10000100;
   // assign rom_data[20998]=8'b00101110;
   // assign rom_data[20999]=8'b10000011;
   // assign rom_data[21000]=8'b00101110;
   // assign rom_data[21001]=8'b10000010;
   // assign rom_data[21002]=8'b00101110;
   // assign rom_data[21003]=8'b10000010;
   // assign rom_data[21004]=8'b00101110;
   // assign rom_data[21005]=8'b10000001;
   // assign rom_data[21006]=8'b00101110;
   // assign rom_data[21007]=8'b01111111;
   // assign rom_data[21008]=8'b00101110;
   // assign rom_data[21009]=8'b01111110;
   // assign rom_data[21010]=8'b00101110;
   // assign rom_data[21011]=8'b01111101;
   // assign rom_data[21012]=8'b00101110;
   // assign rom_data[21013]=8'b01111100;
   // assign rom_data[21014]=8'b00101110;
   // assign rom_data[21015]=8'b01111011;
   // assign rom_data[21016]=8'b00101110;
   // assign rom_data[21017]=8'b01111010;
   // assign rom_data[21018]=8'b00101110;
   // assign rom_data[21019]=8'b01111001;
   // assign rom_data[21020]=8'b00101110;
   // assign rom_data[21021]=8'b01110111;
   // assign rom_data[21022]=8'b00101110;
   // assign rom_data[21023]=8'b01110110;
   // assign rom_data[21024]=8'b00101110;
   // assign rom_data[21025]=8'b01110101;
   // assign rom_data[21026]=8'b00101110;
   // assign rom_data[21027]=8'b01110100;
   // assign rom_data[21028]=8'b00101110;
   // assign rom_data[21029]=8'b01110010;
   // assign rom_data[21030]=8'b00101110;
   // assign rom_data[21031]=8'b01110001;
   // assign rom_data[21032]=8'b00101110;
   // assign rom_data[21033]=8'b01110000;
   // assign rom_data[21034]=8'b00101110;
   // assign rom_data[21035]=8'b01101110;
   // assign rom_data[21036]=8'b00101110;
   // assign rom_data[21037]=8'b01101101;
   // assign rom_data[21038]=8'b00101110;
   // assign rom_data[21039]=8'b01101100;
   // assign rom_data[21040]=8'b00101110;
   // assign rom_data[21041]=8'b01101010;
   // assign rom_data[21042]=8'b00101110;
   // assign rom_data[21043]=8'b01101001;
   // assign rom_data[21044]=8'b00101110;
   // assign rom_data[21045]=8'b01100111;
   // assign rom_data[21046]=8'b00101110;
   // assign rom_data[21047]=8'b01100110;
   // assign rom_data[21048]=8'b00101110;
   // assign rom_data[21049]=8'b01100101;
   // assign rom_data[21050]=8'b00101110;
   // assign rom_data[21051]=8'b01100011;
   // assign rom_data[21052]=8'b00101110;
   // assign rom_data[21053]=8'b01100010;
   // assign rom_data[21054]=8'b00101110;
   // assign rom_data[21055]=8'b01100000;
   // assign rom_data[21056]=8'b00101110;
   // assign rom_data[21057]=8'b01011111;
   // assign rom_data[21058]=8'b00101110;
   // assign rom_data[21059]=8'b01011110;
   // assign rom_data[21060]=8'b00101110;
   // assign rom_data[21061]=8'b01011100;
   // assign rom_data[21062]=8'b00101110;
   // assign rom_data[21063]=8'b01011011;
   // assign rom_data[21064]=8'b00101110;
   // assign rom_data[21065]=8'b01011001;
   // assign rom_data[21066]=8'b00101110;
   // assign rom_data[21067]=8'b01011000;
   // assign rom_data[21068]=8'b00101110;
   // assign rom_data[21069]=8'b01010111;
   // assign rom_data[21070]=8'b00101110;
   // assign rom_data[21071]=8'b01010101;
   // assign rom_data[21072]=8'b00101110;
   // assign rom_data[21073]=8'b01010100;
   // assign rom_data[21074]=8'b00101110;
   // assign rom_data[21075]=8'b01010010;
   // assign rom_data[21076]=8'b00101110;
   // assign rom_data[21077]=8'b01010001;
   // assign rom_data[21078]=8'b00101101;
   // assign rom_data[21079]=8'b01010000;
   // assign rom_data[21080]=8'b00101101;
   // assign rom_data[21081]=8'b01001110;
   // assign rom_data[21082]=8'b00101101;
   // assign rom_data[21083]=8'b01001101;
   // assign rom_data[21084]=8'b00101101;
   // assign rom_data[21085]=8'b01001011;
   // assign rom_data[21086]=8'b00101101;
   // assign rom_data[21087]=8'b01001010;
   // assign rom_data[21088]=8'b00101101;
   // assign rom_data[21089]=8'b01001001;
   // assign rom_data[21090]=8'b00101101;
   // assign rom_data[21091]=8'b01000111;
   // assign rom_data[21092]=8'b00101101;
   // assign rom_data[21093]=8'b01000110;
   // assign rom_data[21094]=8'b00101101;
   // assign rom_data[21095]=8'b01000101;
   // assign rom_data[21096]=8'b00101101;
   // assign rom_data[21097]=8'b01000011;
   // assign rom_data[21098]=8'b00101101;
   // assign rom_data[21099]=8'b01000010;
   // assign rom_data[21100]=8'b00101101;
   // assign rom_data[21101]=8'b01000001;
   // assign rom_data[21102]=8'b00101101;
   // assign rom_data[21103]=8'b01000000;
   // assign rom_data[21104]=8'b00101101;
   // assign rom_data[21105]=8'b00111110;
   // assign rom_data[21106]=8'b00101101;
   // assign rom_data[21107]=8'b00111101;
   // assign rom_data[21108]=8'b00101101;
   // assign rom_data[21109]=8'b00111100;
   // assign rom_data[21110]=8'b00101101;
   // assign rom_data[21111]=8'b00111011;
   // assign rom_data[21112]=8'b00101101;
   // assign rom_data[21113]=8'b00111010;
   // assign rom_data[21114]=8'b00101101;
   // assign rom_data[21115]=8'b00111001;
   // assign rom_data[21116]=8'b00101101;
   // assign rom_data[21117]=8'b00110111;
   // assign rom_data[21118]=8'b00101101;
   // assign rom_data[21119]=8'b00110110;
   // assign rom_data[21120]=8'b00101101;
   // assign rom_data[21121]=8'b00110101;
   // assign rom_data[21122]=8'b00101101;
   // assign rom_data[21123]=8'b00110100;
   // assign rom_data[21124]=8'b00101101;
   // assign rom_data[21125]=8'b00110011;
   // assign rom_data[21126]=8'b00101101;
   // assign rom_data[21127]=8'b00110010;
   // assign rom_data[21128]=8'b00101101;
   // assign rom_data[21129]=8'b00110010;
   // assign rom_data[21130]=8'b00101101;
   // assign rom_data[21131]=8'b00110001;
   // assign rom_data[21132]=8'b00101101;
   // assign rom_data[21133]=8'b00110000;
   // assign rom_data[21134]=8'b00101101;
   // assign rom_data[21135]=8'b00101111;
   // assign rom_data[21136]=8'b00101101;
   // assign rom_data[21137]=8'b00101111;
   // assign rom_data[21138]=8'b00101101;
   // assign rom_data[21139]=8'b00101110;
   // assign rom_data[21140]=8'b00101101;
   // assign rom_data[21141]=8'b00101110;
   // assign rom_data[21142]=8'b00101101;
   // assign rom_data[21143]=8'b00101101;
   // assign rom_data[21144]=8'b00101101;
   // assign rom_data[21145]=8'b00101101;
   // assign rom_data[21146]=8'b00101101;
   // assign rom_data[21147]=8'b00101100;
   // assign rom_data[21148]=8'b00101101;
   // assign rom_data[21149]=8'b00101100;
   // assign rom_data[21150]=8'b00101101;
   // assign rom_data[21151]=8'b00101100;
   // assign rom_data[21152]=8'b00101101;
   // assign rom_data[21153]=8'b00101100;
   // assign rom_data[21154]=8'b00101101;
   // assign rom_data[21155]=8'b00101100;
   // assign rom_data[21156]=8'b00101101;
   // assign rom_data[21157]=8'b00101100;
   // assign rom_data[21158]=8'b00101101;
   // assign rom_data[21159]=8'b00101100;
   // assign rom_data[21160]=8'b00101101;
   // assign rom_data[21161]=8'b00101101;
   // assign rom_data[21162]=8'b00101101;
   // assign rom_data[21163]=8'b00101101;
   // assign rom_data[21164]=8'b00101101;
   // assign rom_data[21165]=8'b00101101;
   // assign rom_data[21166]=8'b00101101;
   // assign rom_data[21167]=8'b00101110;
   // assign rom_data[21168]=8'b00101101;
   // assign rom_data[21169]=8'b00101111;
   // assign rom_data[21170]=8'b00101101;
   // assign rom_data[21171]=8'b00101111;
   // assign rom_data[21172]=8'b00101101;
   // assign rom_data[21173]=8'b00110000;
   // assign rom_data[21174]=8'b00101101;
   // assign rom_data[21175]=8'b00110001;
   // assign rom_data[21176]=8'b00101101;
   // assign rom_data[21177]=8'b00110010;
   // assign rom_data[21178]=8'b00101101;
   // assign rom_data[21179]=8'b00110010;
   // assign rom_data[21180]=8'b00101101;
   // assign rom_data[21181]=8'b00110011;
   // assign rom_data[21182]=8'b00101101;
   // assign rom_data[21183]=8'b00110100;
   // assign rom_data[21184]=8'b00101101;
   // assign rom_data[21185]=8'b00110101;
   // assign rom_data[21186]=8'b00101100;
   // assign rom_data[21187]=8'b00110110;
   // assign rom_data[21188]=8'b00101100;
   // assign rom_data[21189]=8'b00110111;
   // assign rom_data[21190]=8'b00101100;
   // assign rom_data[21191]=8'b00111001;
   // assign rom_data[21192]=8'b00101100;
   // assign rom_data[21193]=8'b00111010;
   // assign rom_data[21194]=8'b00101100;
   // assign rom_data[21195]=8'b00111011;
   // assign rom_data[21196]=8'b00101100;
   // assign rom_data[21197]=8'b00111100;
   // assign rom_data[21198]=8'b00101100;
   // assign rom_data[21199]=8'b00111101;
   // assign rom_data[21200]=8'b00101100;
   // assign rom_data[21201]=8'b00111110;
   // assign rom_data[21202]=8'b00101100;
   // assign rom_data[21203]=8'b01000000;
   // assign rom_data[21204]=8'b00101100;
   // assign rom_data[21205]=8'b01000001;
   // assign rom_data[21206]=8'b00101100;
   // assign rom_data[21207]=8'b01000010;
   // assign rom_data[21208]=8'b00101100;
   // assign rom_data[21209]=8'b01000100;
   // assign rom_data[21210]=8'b00101100;
   // assign rom_data[21211]=8'b01000101;
   // assign rom_data[21212]=8'b00101100;
   // assign rom_data[21213]=8'b01000110;
   // assign rom_data[21214]=8'b00101100;
   // assign rom_data[21215]=8'b01001000;
   // assign rom_data[21216]=8'b00101100;
   // assign rom_data[21217]=8'b01001001;
   // assign rom_data[21218]=8'b00101100;
   // assign rom_data[21219]=8'b01001010;
   // assign rom_data[21220]=8'b00101100;
   // assign rom_data[21221]=8'b01001100;
   // assign rom_data[21222]=8'b00101100;
   // assign rom_data[21223]=8'b01001101;
   // assign rom_data[21224]=8'b00101100;
   // assign rom_data[21225]=8'b01001110;
   // assign rom_data[21226]=8'b00101100;
   // assign rom_data[21227]=8'b01010000;
   // assign rom_data[21228]=8'b00101100;
   // assign rom_data[21229]=8'b01010001;
   // assign rom_data[21230]=8'b00101100;
   // assign rom_data[21231]=8'b01010011;
   // assign rom_data[21232]=8'b00101100;
   // assign rom_data[21233]=8'b01010100;
   // assign rom_data[21234]=8'b00101100;
   // assign rom_data[21235]=8'b01010101;
   // assign rom_data[21236]=8'b00101100;
   // assign rom_data[21237]=8'b01010111;
   // assign rom_data[21238]=8'b00101100;
   // assign rom_data[21239]=8'b01011000;
   // assign rom_data[21240]=8'b00101100;
   // assign rom_data[21241]=8'b01011010;



// reg [23:0] f1_data_d, f1_data_q;
// wire[13:0] f1_addrs;
// reg [15:0] f1_antidata;

reg [23:0] f2_data_d, f2_data_q;
wire[13:0] f2_addrs;
reg [15:0] f2_antidata;

// reg [23:0] f3_data_d, f3_data_q;
// wire[13:0] f3_addrs;
// reg [15:0] f3_antidata;

// reg [23:0] f4_data_d, f4_data_q;
// wire[13:0] f4_addrs;
// reg [15:0] f4_antidata;

// reg [23:0] f5_data_d, f5_data_q;
// wire[13:0] f5_addrs;
// reg [15:0] f5_antidata;

// reg [23:0] f6_data_d, f6_data_q;
// wire[13:0] f6_addrs;
// reg [15:0] f6_antidata;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;

// reg [15:0] f1_CH_A_d, f1_CH_A_q;
// reg [15:0] f1_CH_B_d, f1_CH_B_q;
// reg [15:0] f1_CH_C_d, f1_CH_C_q;
// reg [15:0] f1_CH_D_d, f1_CH_D_q;

reg [15:0] f2_CH_A_d, f2_CH_A_q;
reg [15:0] f2_CH_B_d, f2_CH_B_q;
reg [15:0] f2_CH_C_d, f2_CH_C_q;
reg [15:0] f2_CH_D_d, f2_CH_D_q;

// reg [15:0] f3_CH_A_d, f3_CH_A_q;
// reg [15:0] f3_CH_B_d, f3_CH_B_q;
// reg [15:0] f3_CH_C_d, f3_CH_C_q;
// reg [15:0] f3_CH_D_d, f3_CH_D_q;

// reg [15:0] f4_CH_A_d, f4_CH_A_q;
// reg [15:0] f4_CH_B_d, f4_CH_B_q;
// reg [15:0] f4_CH_C_d, f4_CH_C_q;
// reg [15:0] f4_CH_D_d, f4_CH_D_q;

// reg [15:0] f5_CH_A_d, f5_CH_A_q;
// reg [15:0] f5_CH_B_d, f5_CH_B_q;
// reg [15:0] f5_CH_C_d, f5_CH_C_q;
// reg [15:0] f5_CH_D_d, f5_CH_D_q;

// reg [15:0] f6_CH_A_d, f6_CH_A_q;
// reg [15:0] f6_CH_B_d, f6_CH_B_q;
// reg [15:0] f6_CH_C_d, f6_CH_C_q;
// reg [15:0] f6_CH_D_d, f6_CH_D_q;

// assign f1_data = f1_data_q;
assign f2_data = f2_data_q;
// assign f3_data = f3_data_q;
// assign f4_data = f4_data_q;
// assign f5_data = f5_data_q;
// assign f6_data = f6_data_q;

// assign f1_addrs = f1_addr[15:2];
assign f2_addrs = f2_addr[15:2];
// assign f3_addrs = f3_addr[15:2];
// assign f4_addrs = f4_addr[15:2];
// assign f5_addrs = f5_addr[15:2];
// assign f6_addrs = f6_addr[15:2];

always @(*) begin
    // f1_CH_A_d=f1_CH_A_q;
    // f1_CH_B_d=f1_CH_B_q;
    // f1_CH_C_d=f1_CH_C_q;
    // f1_CH_D_d=f1_CH_D_q;

    f2_CH_A_d=f2_CH_A_q;
    f2_CH_B_d=f2_CH_B_q;
    f2_CH_C_d=f2_CH_C_q;
    f2_CH_D_d=f2_CH_D_q;
    
    // f3_CH_A_d=f3_CH_A_q;
    // f3_CH_B_d=f3_CH_B_q;
    // f3_CH_C_d=f3_CH_C_q;
    // f3_CH_D_d=f3_CH_D_q;
    
    // f4_CH_A_d=f4_CH_A_q;
    // f4_CH_B_d=f4_CH_B_q;
    // f4_CH_C_d=f4_CH_C_q;
    // f4_CH_D_d=f4_CH_D_q;
    
    // f5_CH_A_d=f5_CH_A_q;
    // f5_CH_B_d=f5_CH_B_q;
    // f5_CH_C_d=f5_CH_C_q;
    // f5_CH_D_d=f5_CH_D_q;
    
    // f6_CH_A_d=f6_CH_A_q;
    // f6_CH_B_d=f6_CH_B_q;
    // f6_CH_C_d=f6_CH_C_q;
    // f6_CH_D_d=f6_CH_D_q;


    if (go_home==1'b1) begin
        // F1
        // case (f1_addr[2:1])
        //     2'b00: begin // this is a CHANNEL A
        //         if (f1_CH_A_q>home_bias) begin
        //             f1_CH_A_d=f1_CH_A_q-home_step;
        //         end else if (f1_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f1_CH_A_d=f1_CH_A_q+home_step; 
        //         end 
        //     end
        //     2'b01: begin // this is a CHANNEL C
        //         if (f1_CH_C_q>home_bias) begin
        //             f1_CH_C_d=f1_CH_C_q-home_step;
        //         end else if (f1_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f1_CH_C_d=f1_CH_C_q+home_step;
        //         end 
        //     end
        //     2'b10: begin // this is a CHANNEL B
        //         if (f1_CH_B_q>home_bias) begin
        //             f1_CH_B_d=f1_CH_B_q-home_step;
        //         end else if (f1_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f1_CH_B_d=f1_CH_B_q+home_step; 
        //         end 
        //     end
        //     2'b11: begin // this is a CHANNEL D
        //         if (f1_CH_D_q>home_bias) begin
        //             f1_CH_D_d=f1_CH_D_q-home_step;
        //         end else if (f1_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f1_CH_D_d=f1_CH_D_q+home_step; 
        //         end 
        //     end
        //     default: begin
        //     end
        // endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f2_CH_A_q>home_bias) begin
                    f2_CH_A_d=f2_CH_A_q-home_step;
                end else if (f2_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_A_d=f2_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f2_CH_C_q>home_bias) begin
                    f2_CH_C_d=f2_CH_C_q-home_step;
                end else if (f2_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_C_d=f2_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f2_CH_B_q>home_bias) begin
                    f2_CH_B_d=f2_CH_B_q-home_step;
                end else if (f2_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_B_d=f2_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f2_CH_D_q>home_bias) begin
                    f2_CH_D_d=f2_CH_D_q-home_step;
                end else if (f2_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_D_d=f2_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // // F3
        // case (f3_addr[2:1])
        //     2'b00: begin // this is a CHANNEL A
        //         if (f3_CH_A_q>home_bias) begin
        //             f3_CH_A_d=f3_CH_A_q-home_step;
        //         end else if (f3_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f3_CH_A_d=f3_CH_A_q+home_step; 
        //         end 
        //     end
        //     2'b01: begin // this is a CHANNEL C
        //         if (f3_CH_C_q>home_bias) begin
        //             f3_CH_C_d=f3_CH_C_q-home_step;
        //         end else if (f3_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f3_CH_C_d=f3_CH_C_q+home_step;
        //         end 
        //     end
        //     2'b10: begin // this is a CHANNEL B
        //         if (f3_CH_B_q>home_bias) begin
        //             f3_CH_B_d=f3_CH_B_q-home_step;
        //         end else if (f3_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f3_CH_B_d=f3_CH_B_q+home_step; 
        //         end 
        //     end
        //     2'b11: begin // this is a CHANNEL D
        //         if (f3_CH_D_q>home_bias) begin
        //             f3_CH_D_d=f3_CH_D_q-home_step;
        //         end else if (f3_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f3_CH_D_d=f3_CH_D_q+home_step; 
        //         end 
        //     end
        //     default: begin
        //     end
        // endcase
        // // F4
        // case (f4_addr[2:1])
        //     2'b00: begin // this is a CHANNEL A
        //         if (f4_CH_A_q>home_bias) begin
        //             f4_CH_A_d=f4_CH_A_q-home_step;
        //         end else if (f4_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f4_CH_A_d=f4_CH_A_q+home_step; 
        //         end 
        //     end
        //     2'b01: begin // this is a CHANNEL C
        //         if (f4_CH_C_q>home_bias) begin
        //             f4_CH_C_d=f4_CH_C_q-home_step;
        //         end else if (f4_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f4_CH_C_d=f4_CH_C_q+home_step;
        //         end 
        //     end
        //     2'b10: begin // this is a CHANNEL B
        //         if (f4_CH_B_q>home_bias) begin
        //             f4_CH_B_d=f4_CH_B_q-home_step;
        //         end else if (f4_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f4_CH_B_d=f4_CH_B_q+home_step; 
        //         end 
        //     end
        //     2'b11: begin // this is a CHANNEL D
        //         if (f4_CH_D_q>home_bias) begin
        //             f4_CH_D_d=f4_CH_D_q-home_step;
        //         end else if (f4_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f4_CH_D_d=f4_CH_D_q+home_step; 
        //         end 
        //     end
        //     default: begin
        //     end
        // endcase
        // // F5
        // case (f5_addr[2:1])
        //     2'b00: begin // this is a CHANNEL A
        //         if (f5_CH_A_q>home_bias) begin
        //             f5_CH_A_d=f5_CH_A_q-home_step;
        //         end else if (f5_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f5_CH_A_d=f5_CH_A_q+home_step; 
        //         end 
        //     end
        //     2'b01: begin // this is a CHANNEL C
        //         if (f5_CH_C_q>home_bias) begin
        //             f5_CH_C_d=f5_CH_C_q-home_step;
        //         end else if (f5_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f5_CH_C_d=f5_CH_C_q+home_step;
        //         end 
        //     end
        //     2'b10: begin // this is a CHANNEL B
        //         if (f5_CH_B_q>home_bias) begin
        //             f5_CH_B_d=f5_CH_B_q-home_step;
        //         end else if (f5_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f5_CH_B_d=f5_CH_B_q+home_step; 
        //         end 
        //     end
        //     2'b11: begin // this is a CHANNEL D
        //         if (f5_CH_D_q>home_bias) begin
        //             f5_CH_D_d=f5_CH_D_q-home_step;
        //         end else if (f5_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f5_CH_D_d=f5_CH_D_q+home_step; 
        //         end 
        //     end
        //     default: begin
        //     end
        // endcase
        // // F6
        // case (f6_addr[2:1])
        //     2'b00: begin // this is a CHANNEL A
        //         if (f6_CH_A_q>home_bias) begin
        //             f6_CH_A_d=f6_CH_A_q-home_step;
        //         end else if (f6_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f6_CH_A_d=f6_CH_A_q+home_step; 
        //         end 
        //     end
        //     2'b01: begin // this is a CHANNEL C
        //         if (f6_CH_C_q>home_bias) begin
        //             f6_CH_C_d=f6_CH_C_q-home_step;
        //         end else if (f6_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f6_CH_C_d=f6_CH_C_q+home_step;
        //         end 
        //     end
        //     2'b10: begin // this is a CHANNEL B
        //         if (f6_CH_B_q>home_bias) begin
        //             f6_CH_B_d=f6_CH_B_q-home_step;
        //         end else if (f6_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f6_CH_B_d=f6_CH_B_q+home_step; 
        //         end 
        //     end
        //     2'b11: begin // this is a CHANNEL D
        //         if (f6_CH_D_q>home_bias) begin
        //             f6_CH_D_d=f6_CH_D_q-home_step;
        //         end else if (f6_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
        //             f6_CH_D_d=f6_CH_D_q+home_step; 
        //         end 
        //     end
        //     default: begin
        //     end
        // endcase
    end else begin // if NOT go home
        // // F1
        // case (f1_addr[2:1])
        //     2'b00: begin
        //         f1_CH_A_d= {rom_data[f1_addrs], 8'b10000000};
        //     end
        //     2'b01: begin
        //         f1_CH_C_d= {f1_antidata, 8'b10000000};
        //     end
        //     2'b10: begin
        //         f1_CH_B_d= {rom_data[f1_addrs], 8'b10000000};
        //     end
        //     2'b11: begin
        //         f1_CH_D_d= {f1_antidata, 8'b10000000};
        //     end
        // default: begin
        //     end
        // endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin
                f2_CH_A_d= {rom_data[f2_addrs], 8'b10000000};
            end
            2'b01: begin
                f2_CH_C_d= {f2_antidata, 8'b10000000};
            end
            2'b10: begin
                f2_CH_B_d= {rom_data[f2_addrs],8'b10000000};
            end
            2'b11: begin
                f2_CH_D_d= {f2_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // // F3
        // case (f3_addr[2:1])
        //     2'b00: begin
        //         f3_CH_A_d= {rom_data[f3_addrs], 8'b10000000};
        //     end
        //     2'b01: begin
        //         f3_CH_C_d= {f3_antidata, 8'b10000000};
        //     end
        //     2'b10: begin
        //         f3_CH_B_d= {rom_data[f3_addrs], 8'b10000000};
        //     end
        //     2'b11: begin
        //         f3_CH_D_d= {f3_antidata, 8'b10000000};
        //     end
        // default: begin
        //     end
        // endcase
        // // F4
        // case (f4_addr[2:1])
        //     2'b00: begin
        //         f4_CH_A_d= {rom_data[f4_addrs],8'b10000000};
        //     end
        //     2'b01: begin
        //         f4_CH_C_d= {f4_antidata, 8'b10000000};
        //     end
        //     2'b10: begin
        //         f4_CH_B_d= {rom_data[f4_addrs],8'b10000000};
        //     end
        //     2'b11: begin
        //         f4_CH_D_d= {f4_antidata, 8'b10000000};
        //     end
        // default: begin
        //     end
        // endcase
        // // F5
        // case (f5_addr[2:1])
        //     2'b00: begin
        //         f5_CH_A_d= {rom_data[f5_addrs],8'b10000000};
        //     end
        //     2'b01: begin
        //         f5_CH_C_d= {f5_antidata, 8'b10000000};
        //     end
        //     2'b10: begin
        //         f5_CH_B_d= {rom_data[f5_addrs],8'b10000000};
        //     end
        //     2'b11: begin
        //         f5_CH_D_d= {f5_antidata, 8'b10000000};
        //     end
        // default: begin
        //     end
        // endcase
        // // F6
        // case (f6_addr[2:1])
        //     2'b00: begin
        //         f6_CH_A_d= {rom_data[f6_addrs],8'b10000000};
        //     end
        //     2'b01: begin
        //         f6_CH_C_d= {f6_antidata, 8'b10000000};
        //     end
        //     2'b10: begin
        //         f6_CH_B_d= {rom_data[f6_addrs],8'b10000000};
        //     end
        //     2'b11: begin
        //         f6_CH_D_d= {f6_antidata, 8'b10000000};
        //     end
        // default: begin
        //     end
        // endcase

    end // if go home 

end // always

always @(*) begin
  // f1_antidata = 8'hB4 - rom_data[f1_addrs];
  f2_antidata = 8'hB4 - rom_data[f2_addrs];
  // f3_antidata = 8'hB4 - rom_data[f3_addrs];
  // f4_antidata = 8'hB4 - rom_data[f4_addrs];
  // f5_antidata = 8'hB4 - rom_data[f5_addrs];
  // f6_antidata = 8'hB4 - rom_data[f6_addrs];

 
  // // F1   
  // if (f1_addr==0) begin
  //   f1_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  // end else if (f1_addr==1) begin
  //   f1_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  // end else if (f1_addr[0]==1'b0) begin
  //   f1_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  // end else begin //data in 50%
  //       case (f1_addr[2:1])
  //           2'b00: begin // this is a CHANNEL A
  //               f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_A_q};
  //           end
  //           2'b01: begin // this is a CHANNEL C
  //               f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_C_q};
  //           end
  //           2'b10: begin // this is a CHANNEL B
  //               f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_B_q};
  //           end
  //           2'b11: begin // this is a CHANNEL D
  //               f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_D_q};
  //           end
  //           default: begin
  //           end
  //       endcase
  //  end // if addr=0
  // F2
  if (f2_addr==0) begin
    f2_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f2_addr==1) begin
    f2_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f2_addr[0]==1'b0) begin
    f2_data_d = 24'b00111000_0000000000000000; // Vref send in 50% samples  
  end else begin //data in 50%
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_D_q};
            end
            default: begin
            end
        endcase
   end // if addr=0
  // // F3
  // if (f3_addr==0) begin
  //   f3_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  // end else if (f3_addr==1) begin
  //   f3_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  // end else if (f3_addr[0]==1'b0) begin
  //   f3_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  // end else begin //data in 50%
  //       case (f3_addr[2:1])
  //           2'b00: begin // this is a CHANNEL A
  //               f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_A_q};
  //           end
  //           2'b01: begin // this is a CHANNEL C
  //               f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_C_q};
  //           end
  //           2'b10: begin // this is a CHANNEL B
  //               f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_B_q};
  //           end
  //           2'b11: begin // this is a CHANNEL D
  //               f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_D_q};
  //           end
  //           default: begin
  //           end
  //       endcase
  // end // if addr=0
  // // F4
  // if (f4_addr==0) begin
  //   f4_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  // end else if (f4_addr==1) begin
  //   f4_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  // end else if (f4_addr[0]==1'b0) begin
  //   f4_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  // end else begin //data in 50%
  //       case (f4_addr[2:1])
  //           2'b00: begin // this is a CHANNEL A
  //               f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_A_q};
  //           end
  //           2'b01: begin // this is a CHANNEL C
  //               f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_C_q};
  //           end
  //           2'b10: begin // this is a CHANNEL B
  //               f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_B_q};
  //           end
  //           2'b11: begin // this is a CHANNEL D
  //               f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_D_q};
  //           end
  //           default: begin
  //           end
  //       endcase
  // end // if addr=0
  // // F5
  // if (f5_addr==0) begin
  //   f5_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  // end else if (f5_addr==1) begin
  //   f5_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  // end else if (f5_addr[0]==1'b0) begin
  //   f5_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  // end else begin //data in 50%
  //       case (f5_addr[2:1])
  //           2'b00: begin // this is a CHANNEL A
  //               f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_A_q};
  //           end
  //           2'b01: begin // this is a CHANNEL C
  //               f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_C_q};
  //           end
  //           2'b10: begin // this is a CHANNEL B
  //               f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_B_q};
  //           end
  //           2'b11: begin // this is a CHANNEL D
  //               f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_D_q};
  //           end
  //           default: begin
  //           end
  //       endcase
  // end // if addr=0
  // // F6
  // if (f6_addr==0) begin
  //   f6_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  // end else if (f6_addr==1) begin
  //   f6_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  // end else if (f6_addr[0]==1'b0) begin
  //   f6_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  // end else begin //data in 50%
  //       case (f6_addr[2:1])
  //           2'b00: begin // this is a CHANNEL A
  //               f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_A_q};
  //           end
  //           2'b01: begin // this is a CHANNEL C
  //               f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_C_q};
  //           end
  //           2'b10: begin // this is a CHANNEL B
  //               f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_B_q};
  //           end
  //           2'b11: begin // this is a CHANNEL D
  //               f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_D_q};
  //           end
  //           default: begin
  //           end
  //       endcase
  // end // if addr=0
end // always

// always @(posedge f1_addr[0]) begin
//     f1_CH_A_q<=f1_CH_A_d;
//     f1_CH_B_q<=f1_CH_B_d;
//     f1_CH_C_q<=f1_CH_C_d;
//     f1_CH_D_q<=f1_CH_D_d;
// end

always @(posedge f2_addr[0]) begin
    f2_CH_A_q<=f2_CH_A_d;
    f2_CH_B_q<=f2_CH_B_d;
    f2_CH_C_q<=f2_CH_C_d;
    f2_CH_D_q<=f2_CH_D_d;
end

// always @(posedge f3_addr[0]) begin
//     f3_CH_A_q<=f3_CH_A_d;
//     f3_CH_B_q<=f3_CH_B_d;
//     f3_CH_C_q<=f3_CH_C_d;
//     f3_CH_D_q<=f3_CH_D_d;
// end

// always @(posedge f4_addr[0]) begin
//     f4_CH_A_q<=f4_CH_A_d;
//     f4_CH_B_q<=f4_CH_B_d;
//     f4_CH_C_q<=f4_CH_C_d;
//     f4_CH_D_q<=f4_CH_D_d;
// end

// always @(posedge f5_addr[0]) begin
//     f5_CH_A_q<=f5_CH_A_d;
//     f5_CH_B_q<=f5_CH_B_d;
//     f5_CH_C_q<=f5_CH_C_d;
//     f5_CH_D_q<=f5_CH_D_d;
// end

// always @(posedge f6_addr[0]) begin
//     f6_CH_A_q<=f6_CH_A_d;
//     f6_CH_B_q<=f6_CH_B_d;
//     f6_CH_C_q<=f6_CH_C_d;
//     f6_CH_D_q<=f6_CH_D_d;
// end

always @(posedge clk) begin
    // f1_data_q <= f1_data_d;
    f2_data_q <= f2_data_d;
    // f3_data_q <= f3_data_d;
    // f4_data_q <= f4_data_d;
    // f5_data_q <= f5_data_d;
    // f6_data_q <= f6_data_d;
end // always
 
endmodule