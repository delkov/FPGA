module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] f1_addr,
    input [15:0] f2_addr,
    input [15:0] f3_addr,
    input [15:0] f4_addr,
    input [15:0] f5_addr,
    input [15:0] f6_addr,

    input go_home,
    // OUTPUT
    output [23:0] f1_data,
    output [23:0] f2_data,
    output [23:0] f3_data,
    output [23:0] f4_data,
    output [23:0] f5_data,
    output [23:0] f6_data
  );
  
parameter rom_size = 3241;

reg [7:0] rom_data [rom_size:0];

reg [23:0] f1_data_d, f1_data_q;
wire[13:0] f1_addrs;
reg [15:0] f1_antidata;

reg [23:0] f2_data_d, f2_data_q;
wire[13:0] f2_addrs;
reg [15:0] f2_antidata;

reg [23:0] f3_data_d, f3_data_q;
wire[13:0] f3_addrs;
reg [15:0] f3_antidata;

reg [23:0] f4_data_d, f4_data_q;
wire[13:0] f4_addrs;
reg [15:0] f4_antidata;

reg [23:0] f5_data_d, f5_data_q;
wire[13:0] f5_addrs;
reg [15:0] f5_antidata;

reg [23:0] f6_data_d, f6_data_q;
wire[13:0] f6_addrs;
reg [15:0] f6_antidata;

reg done;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;

reg [15:0] f1_CH_A_d, f1_CH_A_q;
reg [15:0] f1_CH_B_d, f1_CH_B_q;
reg [15:0] f1_CH_C_d, f1_CH_C_q;
reg [15:0] f1_CH_D_d, f1_CH_D_q;

reg [15:0] f2_CH_A_d, f2_CH_A_q;
reg [15:0] f2_CH_B_d, f2_CH_B_q;
reg [15:0] f2_CH_C_d, f2_CH_C_q;
reg [15:0] f2_CH_D_d, f2_CH_D_q;

reg [15:0] f3_CH_A_d, f3_CH_A_q;
reg [15:0] f3_CH_B_d, f3_CH_B_q;
reg [15:0] f3_CH_C_d, f3_CH_C_q;
reg [15:0] f3_CH_D_d, f3_CH_D_q;

reg [15:0] f4_CH_A_d, f4_CH_A_q;
reg [15:0] f4_CH_B_d, f4_CH_B_q;
reg [15:0] f4_CH_C_d, f4_CH_C_q;
reg [15:0] f4_CH_D_d, f4_CH_D_q;

reg [15:0] f5_CH_A_d, f5_CH_A_q;
reg [15:0] f5_CH_B_d, f5_CH_B_q;
reg [15:0] f5_CH_C_d, f5_CH_C_q;
reg [15:0] f5_CH_D_d, f5_CH_D_q;

reg [15:0] f6_CH_A_d, f6_CH_A_q;
reg [15:0] f6_CH_B_d, f6_CH_B_q;
reg [15:0] f6_CH_C_d, f6_CH_C_q;
reg [15:0] f6_CH_D_d, f6_CH_D_q;

assign f1_data = f1_data_q;
assign f2_data = f2_data_q;
assign f3_data = f3_data_q;
assign f4_data = f4_data_q;
assign f5_data = f5_data_q;
assign f6_data = f6_data_q;

assign f1_addrs = f1_addr[15:2];
assign f2_addrs = f2_addr[15:2];
assign f3_addrs = f3_addr[15:2];
assign f4_addrs = f4_addr[15:2];
assign f5_addrs = f5_addr[15:2];
assign f6_addrs = f6_addr[15:2];

always @(*) begin
    f1_CH_A_d=f1_CH_A_q;
    f1_CH_B_d=f1_CH_B_q;
    f1_CH_C_d=f1_CH_C_q;
    f1_CH_D_d=f1_CH_D_q;

    f2_CH_A_d=f2_CH_A_q;
    f2_CH_B_d=f2_CH_B_q;
    f2_CH_C_d=f2_CH_C_q;
    f2_CH_D_d=f2_CH_D_q;
    
    f3_CH_A_d=f3_CH_A_q;
    f3_CH_B_d=f3_CH_B_q;
    f3_CH_C_d=f3_CH_C_q;
    f3_CH_D_d=f3_CH_D_q;
    
    f4_CH_A_d=f4_CH_A_q;
    f4_CH_B_d=f4_CH_B_q;
    f4_CH_C_d=f4_CH_C_q;
    f4_CH_D_d=f4_CH_D_q;
    
    f5_CH_A_d=f5_CH_A_q;
    f5_CH_B_d=f5_CH_B_q;
    f5_CH_C_d=f5_CH_C_q;
    f5_CH_D_d=f5_CH_D_q;
    
    f6_CH_A_d=f6_CH_A_q;
    f6_CH_B_d=f6_CH_B_q;
    f6_CH_C_d=f6_CH_C_q;
    f6_CH_D_d=f6_CH_D_q;


    if (go_home==1'b1) begin
        // F1
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f1_CH_A_q>home_bias) begin
                    f1_CH_A_d=f1_CH_A_q-home_step;
                end else if (f1_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_A_d=f1_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f1_CH_C_q>home_bias) begin
                    f1_CH_C_d=f1_CH_C_q-home_step;
                end else if (f1_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_C_d=f1_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f1_CH_B_q>home_bias) begin
                    f1_CH_B_d=f1_CH_B_q-home_step;
                end else if (f1_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_B_d=f1_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f1_CH_D_q>home_bias) begin
                    f1_CH_D_d=f1_CH_D_q-home_step;
                end else if (f1_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_D_d=f1_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f2_CH_A_q>home_bias) begin
                    f2_CH_A_d=f2_CH_A_q-home_step;
                end else if (f2_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_A_d=f2_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f2_CH_C_q>home_bias) begin
                    f2_CH_C_d=f2_CH_C_q-home_step;
                end else if (f2_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_C_d=f2_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f2_CH_B_q>home_bias) begin
                    f2_CH_B_d=f2_CH_B_q-home_step;
                end else if (f2_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_B_d=f2_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f2_CH_D_q>home_bias) begin
                    f2_CH_D_d=f2_CH_D_q-home_step;
                end else if (f2_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_D_d=f2_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F3
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f3_CH_A_q>home_bias) begin
                    f3_CH_A_d=f3_CH_A_q-home_step;
                end else if (f3_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_A_d=f3_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f3_CH_C_q>home_bias) begin
                    f3_CH_C_d=f3_CH_C_q-home_step;
                end else if (f3_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_C_d=f3_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f3_CH_B_q>home_bias) begin
                    f3_CH_B_d=f3_CH_B_q-home_step;
                end else if (f3_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_B_d=f3_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f3_CH_D_q>home_bias) begin
                    f3_CH_D_d=f3_CH_D_q-home_step;
                end else if (f3_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_D_d=f3_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F4
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f4_CH_A_q>home_bias) begin
                    f4_CH_A_d=f4_CH_A_q-home_step;
                end else if (f4_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_A_d=f4_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f4_CH_C_q>home_bias) begin
                    f4_CH_C_d=f4_CH_C_q-home_step;
                end else if (f4_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_C_d=f4_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f4_CH_B_q>home_bias) begin
                    f4_CH_B_d=f4_CH_B_q-home_step;
                end else if (f4_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_B_d=f4_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f4_CH_D_q>home_bias) begin
                    f4_CH_D_d=f4_CH_D_q-home_step;
                end else if (f4_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_D_d=f4_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F5
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f5_CH_A_q>home_bias) begin
                    f5_CH_A_d=f5_CH_A_q-home_step;
                end else if (f5_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_A_d=f5_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f5_CH_C_q>home_bias) begin
                    f5_CH_C_d=f5_CH_C_q-home_step;
                end else if (f5_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_C_d=f5_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f5_CH_B_q>home_bias) begin
                    f5_CH_B_d=f5_CH_B_q-home_step;
                end else if (f5_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_B_d=f5_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f5_CH_D_q>home_bias) begin
                    f5_CH_D_d=f5_CH_D_q-home_step;
                end else if (f5_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_D_d=f5_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F6
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f6_CH_A_q>home_bias) begin
                    f6_CH_A_d=f6_CH_A_q-home_step;
                end else if (f6_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_A_d=f6_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f6_CH_C_q>home_bias) begin
                    f6_CH_C_d=f6_CH_C_q-home_step;
                end else if (f6_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_C_d=f6_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f6_CH_B_q>home_bias) begin
                    f6_CH_B_d=f6_CH_B_q-home_step;
                end else if (f6_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_B_d=f6_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f6_CH_D_q>home_bias) begin
                    f6_CH_D_d=f6_CH_D_q-home_step;
                end else if (f6_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_D_d=f6_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
    end else begin // if NOT go home
        // F1
        case (f1_addr[2:1])
            2'b00: begin
                f1_CH_A_d= {rom_data[f1_addrs], 8'b10000000};
            end
            2'b01: begin
                f1_CH_C_d= {f1_antidata, 8'b10000000};
            end
            2'b10: begin
                f1_CH_B_d= {rom_data[f1_addrs], 8'b10000000};
            end
            2'b11: begin
                f1_CH_D_d= {f1_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin
                f2_CH_A_d= {rom_data[f2_addrs], 8'b10000000};
            end
            2'b01: begin
                f2_CH_C_d= {f2_antidata, 8'b10000000};
            end
            2'b10: begin
                f2_CH_B_d= {rom_data[f2_addrs],8'b10000000};
            end
            2'b11: begin
                f2_CH_D_d= {f2_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F3
        case (f3_addr[2:1])
            2'b00: begin
                f3_CH_A_d= {rom_data[f3_addrs], 8'b10000000};
            end
            2'b01: begin
                f3_CH_C_d= {f3_antidata, 8'b10000000};
            end
            2'b10: begin
                f3_CH_B_d= {rom_data[f3_addrs], 8'b10000000};
            end
            2'b11: begin
                f3_CH_D_d= {f3_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F4
        case (f4_addr[2:1])
            2'b00: begin
                f4_CH_A_d= {rom_data[f4_addrs],8'b10000000};
            end
            2'b01: begin
                f4_CH_C_d= {f4_antidata, 8'b10000000};
            end
            2'b10: begin
                f4_CH_B_d= {rom_data[f4_addrs],8'b10000000};
            end
            2'b11: begin
                f4_CH_D_d= {f4_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F5
        case (f5_addr[2:1])
            2'b00: begin
                f5_CH_A_d= {rom_data[f5_addrs],8'b10000000};
            end
            2'b01: begin
                f5_CH_C_d= {f5_antidata, 8'b10000000};
            end
            2'b10: begin
                f5_CH_B_d= {rom_data[f5_addrs],8'b10000000};
            end
            2'b11: begin
                f5_CH_D_d= {f5_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F6
        case (f6_addr[2:1])
            2'b00: begin
                f6_CH_A_d= {rom_data[f6_addrs],8'b10000000};
            end
            2'b01: begin
                f6_CH_C_d= {f6_antidata, 8'b10000000};
            end
            2'b10: begin
                f6_CH_B_d= {rom_data[f6_addrs],8'b10000000};
            end
            2'b11: begin
                f6_CH_D_d= {f6_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase

    end // if go home 

end // always

always @(*) begin
  f1_antidata = 8'hB4 - rom_data[f1_addrs];
  f2_antidata = 8'hB4 - rom_data[f2_addrs];
  f3_antidata = 8'hB4 - rom_data[f3_addrs];
  f4_antidata = 8'hB4 - rom_data[f4_addrs];
  f5_antidata = 8'hB4 - rom_data[f5_addrs];
  f6_antidata = 8'hB4 - rom_data[f6_addrs];

    rom_data[ 2]=8'b00101101;
    rom_data[ 3]=8'b01011011;
    rom_data[ 4]=8'b00101101;
    rom_data[ 5]=8'b01011100;
    rom_data[ 6]=8'b00101101;
    rom_data[ 7]=8'b01011110;
    rom_data[ 8]=8'b00101101;
    rom_data[ 9]=8'b01011111;
    rom_data[10]=8'b00101101;
    rom_data[11]=8'b01100001;
    rom_data[12]=8'b00101101;
    rom_data[13]=8'b01100010;
    rom_data[14]=8'b00101101;
    rom_data[15]=8'b01100011;
    rom_data[16]=8'b00101101;
    rom_data[17]=8'b01100101;
    rom_data[18]=8'b00101110;
    rom_data[19]=8'b01100110;
    rom_data[20]=8'b00101110;
    rom_data[21]=8'b01100111;
    rom_data[22]=8'b00101110;
    rom_data[23]=8'b01101001;
    rom_data[24]=8'b00101110;
    rom_data[25]=8'b01101010;
    rom_data[26]=8'b00101110;
    rom_data[27]=8'b01101100;
    rom_data[28]=8'b00101110;
    rom_data[29]=8'b01101101;
    rom_data[30]=8'b00101110;
    rom_data[31]=8'b01101110;
    rom_data[32]=8'b00101110;
    rom_data[33]=8'b01110000;
    rom_data[34]=8'b00101110;
    rom_data[35]=8'b01110001;
    rom_data[36]=8'b00101110;
    rom_data[37]=8'b01110010;
    rom_data[38]=8'b00101110;
    rom_data[39]=8'b01110100;
    rom_data[40]=8'b00101110;
    rom_data[41]=8'b01110101;
    rom_data[42]=8'b00101110;
    rom_data[43]=8'b01110110;
    rom_data[44]=8'b00101110;
    rom_data[45]=8'b01110111;
    rom_data[46]=8'b00101111;
    rom_data[47]=8'b01111001;
    rom_data[48]=8'b00101111;
    rom_data[49]=8'b01111010;
    rom_data[50]=8'b00101111;
    rom_data[51]=8'b01111011;
    rom_data[52]=8'b00101111;
    rom_data[53]=8'b01111100;
    rom_data[54]=8'b00101111;
    rom_data[55]=8'b01111101;
    rom_data[56]=8'b00101111;
    rom_data[57]=8'b01111110;
    rom_data[58]=8'b00101111;
    rom_data[59]=8'b01111111;
    rom_data[60]=8'b00101111;
    rom_data[61]=8'b10000000;
    rom_data[62]=8'b00101111;
    rom_data[63]=8'b10000001;
    rom_data[64]=8'b00110000;
    rom_data[65]=8'b10000010;
    rom_data[66]=8'b00110000;
    rom_data[67]=8'b10000011;
    rom_data[68]=8'b00110000;
    rom_data[69]=8'b10000100;
    rom_data[70]=8'b00110000;
    rom_data[71]=8'b10000101;
    rom_data[72]=8'b00110000;
    rom_data[73]=8'b10000110;
    rom_data[74]=8'b00110000;
    rom_data[75]=8'b10000110;
    rom_data[76]=8'b00110000;
    rom_data[77]=8'b10000111;
    rom_data[78]=8'b00110000;
    rom_data[79]=8'b10001000;
    rom_data[80]=8'b00110000;
    rom_data[81]=8'b10001000;
    rom_data[82]=8'b00110001;
    rom_data[83]=8'b10001001;
    rom_data[84]=8'b00110001;
    rom_data[85]=8'b10001001;
    rom_data[86]=8'b00110001;
    rom_data[87]=8'b10001001;
    rom_data[88]=8'b00110001;
    rom_data[89]=8'b10001010;
    rom_data[90]=8'b00110001;
    rom_data[91]=8'b10001010;
    rom_data[92]=8'b00110001;
    rom_data[93]=8'b10001010;
    rom_data[94]=8'b00110001;
    rom_data[95]=8'b10001010;
    rom_data[96]=8'b00110010;
    rom_data[97]=8'b10001010;
    rom_data[98]=8'b00110010;
    rom_data[99]=8'b10001001;
    rom_data[100]=8'b00110010;
    rom_data[101]=8'b10001001;
    rom_data[102]=8'b00110010;
    rom_data[103]=8'b10001001;
    rom_data[104]=8'b00110010;
    rom_data[105]=8'b10001000;
    rom_data[106]=8'b00110010;
    rom_data[107]=8'b10001000;
    rom_data[108]=8'b00110010;
    rom_data[109]=8'b10000111;
    rom_data[110]=8'b00110010;
    rom_data[111]=8'b10000111;
    rom_data[112]=8'b00110011;
    rom_data[113]=8'b10000110;
    rom_data[114]=8'b00110011;
    rom_data[115]=8'b10000101;
    rom_data[116]=8'b00110011;
    rom_data[117]=8'b10000100;
    rom_data[118]=8'b00110011;
    rom_data[119]=8'b10000011;
    rom_data[120]=8'b00110011;
    rom_data[121]=8'b10000011;
    rom_data[122]=8'b00110011;
    rom_data[123]=8'b10000010;
    rom_data[124]=8'b00110011;
    rom_data[125]=8'b10000001;
    rom_data[126]=8'b00110011;
    rom_data[127]=8'b10000000;
    rom_data[128]=8'b00110100;
    rom_data[129]=8'b01111110;
    rom_data[130]=8'b00110100;
    rom_data[131]=8'b01111101;
    rom_data[132]=8'b00110100;
    rom_data[133]=8'b01111100;
    rom_data[134]=8'b00110100;
    rom_data[135]=8'b01111011;
    rom_data[136]=8'b00110100;
    rom_data[137]=8'b01111010;
    rom_data[138]=8'b00110100;
    rom_data[139]=8'b01111001;
    rom_data[140]=8'b00110100;
    rom_data[141]=8'b01110111;
    rom_data[142]=8'b00110100;
    rom_data[143]=8'b01110110;
    rom_data[144]=8'b00110101;
    rom_data[145]=8'b01110101;
    rom_data[146]=8'b00110101;
    rom_data[147]=8'b01110100;
    rom_data[148]=8'b00110101;
    rom_data[149]=8'b01110010;
    rom_data[150]=8'b00110101;
    rom_data[151]=8'b01110001;
    rom_data[152]=8'b00110101;
    rom_data[153]=8'b01110000;
    rom_data[154]=8'b00110101;
    rom_data[155]=8'b01101110;
    rom_data[156]=8'b00110101;
    rom_data[157]=8'b01101101;
    rom_data[158]=8'b00110101;
    rom_data[159]=8'b01101100;
    rom_data[160]=8'b00110101;
    rom_data[161]=8'b01101010;
    rom_data[162]=8'b00110101;
    rom_data[163]=8'b01101001;
    rom_data[164]=8'b00110110;
    rom_data[165]=8'b01101000;
    rom_data[166]=8'b00110110;
    rom_data[167]=8'b01100110;
    rom_data[168]=8'b00110110;
    rom_data[169]=8'b01100101;
    rom_data[170]=8'b00110110;
    rom_data[171]=8'b01100011;
    rom_data[172]=8'b00110110;
    rom_data[173]=8'b01100010;
    rom_data[174]=8'b00110110;
    rom_data[175]=8'b01100001;
    rom_data[176]=8'b00110110;
    rom_data[177]=8'b01011111;
    rom_data[178]=8'b00110110;
    rom_data[179]=8'b01011110;
    rom_data[180]=8'b00110110;
    rom_data[181]=8'b01011100;
    rom_data[182]=8'b00110110;
    rom_data[183]=8'b01011011;
    rom_data[184]=8'b00110111;
    rom_data[185]=8'b01011010;
    rom_data[186]=8'b00110111;
    rom_data[187]=8'b01011000;
    rom_data[188]=8'b00110111;
    rom_data[189]=8'b01010111;
    rom_data[190]=8'b00110111;
    rom_data[191]=8'b01010101;
    rom_data[192]=8'b00110111;
    rom_data[193]=8'b01010100;
    rom_data[194]=8'b00110111;
    rom_data[195]=8'b01010010;
    rom_data[196]=8'b00110111;
    rom_data[197]=8'b01010001;
    rom_data[198]=8'b00110111;
    rom_data[199]=8'b01010000;
    rom_data[200]=8'b00110111;
    rom_data[201]=8'b01001110;
    rom_data[202]=8'b00110111;
    rom_data[203]=8'b01001101;
    rom_data[204]=8'b00111000;
    rom_data[205]=8'b01001100;
    rom_data[206]=8'b00111000;
    rom_data[207]=8'b01001010;
    rom_data[208]=8'b00111000;
    rom_data[209]=8'b01001001;
    rom_data[210]=8'b00111000;
    rom_data[211]=8'b01001000;
    rom_data[212]=8'b00111000;
    rom_data[213]=8'b01000110;
    rom_data[214]=8'b00111000;
    rom_data[215]=8'b01000101;
    rom_data[216]=8'b00111000;
    rom_data[217]=8'b01000100;
    rom_data[218]=8'b00111000;
    rom_data[219]=8'b01000010;
    rom_data[220]=8'b00111000;
    rom_data[221]=8'b01000001;
    rom_data[222]=8'b00111001;
    rom_data[223]=8'b01000000;
    rom_data[224]=8'b00111001;
    rom_data[225]=8'b00111111;
    rom_data[226]=8'b00111001;
    rom_data[227]=8'b00111101;
    rom_data[228]=8'b00111001;
    rom_data[229]=8'b00111100;
    rom_data[230]=8'b00111001;
    rom_data[231]=8'b00111011;
    rom_data[232]=8'b00111001;
    rom_data[233]=8'b00111010;
    rom_data[234]=8'b00111001;
    rom_data[235]=8'b00111001;
    rom_data[236]=8'b00111001;
    rom_data[237]=8'b00111000;
    rom_data[238]=8'b00111001;
    rom_data[239]=8'b00110110;
    rom_data[240]=8'b00111010;
    rom_data[241]=8'b00110101;
    rom_data[242]=8'b00111010;
    rom_data[243]=8'b00110100;
    rom_data[244]=8'b00111010;
    rom_data[245]=8'b00110011;
    rom_data[246]=8'b00111010;
    rom_data[247]=8'b00110011;
    rom_data[248]=8'b00111010;
    rom_data[249]=8'b00110010;
    rom_data[250]=8'b00111010;
    rom_data[251]=8'b00110001;
    rom_data[252]=8'b00111010;
    rom_data[253]=8'b00110000;
    rom_data[254]=8'b00111010;
    rom_data[255]=8'b00101111;
    rom_data[256]=8'b00111011;
    rom_data[257]=8'b00101111;
    rom_data[258]=8'b00111011;
    rom_data[259]=8'b00101110;
    rom_data[260]=8'b00111011;
    rom_data[261]=8'b00101110;
    rom_data[262]=8'b00111011;
    rom_data[263]=8'b00101101;
    rom_data[264]=8'b00111011;
    rom_data[265]=8'b00101101;
    rom_data[266]=8'b00111011;
    rom_data[267]=8'b00101100;
    rom_data[268]=8'b00111011;
    rom_data[269]=8'b00101100;
    rom_data[270]=8'b00111100;
    rom_data[271]=8'b00101100;
    rom_data[272]=8'b00111100;
    rom_data[273]=8'b00101100;
    rom_data[274]=8'b00111100;
    rom_data[275]=8'b00101100;
    rom_data[276]=8'b00111100;
    rom_data[277]=8'b00101100;
    rom_data[278]=8'b00111100;
    rom_data[279]=8'b00101100;
    rom_data[280]=8'b00111100;
    rom_data[281]=8'b00101101;
    rom_data[282]=8'b00111100;
    rom_data[283]=8'b00101101;
    rom_data[284]=8'b00111100;
    rom_data[285]=8'b00101101;
    rom_data[286]=8'b00111101;
    rom_data[287]=8'b00101110;
    rom_data[288]=8'b00111101;
    rom_data[289]=8'b00101111;
    rom_data[290]=8'b00111101;
    rom_data[291]=8'b00101111;
    rom_data[292]=8'b00111101;
    rom_data[293]=8'b00110000;
    rom_data[294]=8'b00111101;
    rom_data[295]=8'b00110001;
    rom_data[296]=8'b00111101;
    rom_data[297]=8'b00110001;
    rom_data[298]=8'b00111101;
    rom_data[299]=8'b00110010;
    rom_data[300]=8'b00111110;
    rom_data[301]=8'b00110011;
    rom_data[302]=8'b00111110;
    rom_data[303]=8'b00110100;
    rom_data[304]=8'b00111110;
    rom_data[305]=8'b00110101;
    rom_data[306]=8'b00111110;
    rom_data[307]=8'b00110110;
    rom_data[308]=8'b00111110;
    rom_data[309]=8'b00110111;
    rom_data[310]=8'b00111110;
    rom_data[311]=8'b00111000;
    rom_data[312]=8'b00111110;
    rom_data[313]=8'b00111010;
    rom_data[314]=8'b00111110;
    rom_data[315]=8'b00111011;
    rom_data[316]=8'b00111110;
    rom_data[317]=8'b00111100;
    rom_data[318]=8'b00111111;
    rom_data[319]=8'b00111101;
    rom_data[320]=8'b00111111;
    rom_data[321]=8'b00111110;
    rom_data[322]=8'b00111111;
    rom_data[323]=8'b01000000;
    rom_data[324]=8'b00111111;
    rom_data[325]=8'b01000001;
    rom_data[326]=8'b00111111;
    rom_data[327]=8'b01000010;
    rom_data[328]=8'b00111111;
    rom_data[329]=8'b01000100;
    rom_data[330]=8'b00111111;
    rom_data[331]=8'b01000101;
    rom_data[332]=8'b00111111;
    rom_data[333]=8'b01000110;
    rom_data[334]=8'b00111111;
    rom_data[335]=8'b01000111;
    rom_data[336]=8'b01000000;
    rom_data[337]=8'b01001001;
    rom_data[338]=8'b01000000;
    rom_data[339]=8'b01001010;
    rom_data[340]=8'b01000000;
    rom_data[341]=8'b01001100;
    rom_data[342]=8'b01000000;
    rom_data[343]=8'b01001101;
    rom_data[344]=8'b01000000;
    rom_data[345]=8'b01001110;
    rom_data[346]=8'b01000000;
    rom_data[347]=8'b01010000;
    rom_data[348]=8'b01000000;
    rom_data[349]=8'b01010001;
    rom_data[350]=8'b01000000;
    rom_data[351]=8'b01010010;
    rom_data[352]=8'b01000000;
    rom_data[353]=8'b01010100;
    rom_data[354]=8'b01000000;
    rom_data[355]=8'b01010101;
    rom_data[356]=8'b01000001;
    rom_data[357]=8'b01010111;
    rom_data[358]=8'b01000001;
    rom_data[359]=8'b01011000;
    rom_data[360]=8'b01000001;
    rom_data[361]=rom_data[12];
    rom_data[362]=8'b01000001;
    rom_data[363]=rom_data[12];
    rom_data[364]=8'b01000001;
    rom_data[365]=rom_data[12];
    rom_data[366]=8'b01000001;
    rom_data[367]=rom_data[12];
    rom_data[368]=8'b01000001;
    rom_data[369]=rom_data[12];
    rom_data[370]=8'b01000001;
    rom_data[371]=rom_data[12];
    rom_data[372]=8'b01000001;
    rom_data[373]=rom_data[12];
    rom_data[374]=8'b01000001;
    rom_data[375]=rom_data[12];
    rom_data[376]=8'b01000010;
    rom_data[377]=rom_data[12];
    rom_data[378]=8'b01000010;
    rom_data[379]=rom_data[12];
    rom_data[380]=8'b01000010;
    rom_data[381]=rom_data[12];
    rom_data[382]=8'b01000010;
    rom_data[383]=rom_data[12];
    rom_data[384]=8'b01000010;
    rom_data[385]=rom_data[12];
    rom_data[386]=8'b01000010;
    rom_data[387]=rom_data[12];
    rom_data[388]=8'b01000010;
    rom_data[389]=rom_data[12];
    rom_data[390]=8'b01000010;
    rom_data[391]=rom_data[12];
    rom_data[392]=8'b01000010;
    rom_data[393]=rom_data[12];
    rom_data[394]=8'b01000011;
    rom_data[395]=rom_data[12];
    rom_data[396]=8'b01000011;
    rom_data[397]=rom_data[12];
    rom_data[398]=8'b01000011;
    rom_data[399]=rom_data[12];
    rom_data[400]=8'b01000011;
    rom_data[401]=rom_data[12];
    rom_data[402]=8'b01000011;
    rom_data[403]=rom_data[12];
    rom_data[404]=8'b01000011;
    rom_data[405]=rom_data[12];
    rom_data[406]=8'b01000011;
    rom_data[407]=rom_data[12];
    rom_data[408]=8'b01000011;
    rom_data[409]=rom_data[12];
    rom_data[410]=8'b01000011;
    rom_data[411]=rom_data[12];
    rom_data[412]=8'b01000011;
    rom_data[413]=rom_data[12];
    rom_data[414]=8'b01000100;
    rom_data[415]=rom_data[12];
    rom_data[416]=8'b01000100;
    rom_data[417]=rom_data[12];
    rom_data[418]=8'b01000100;
    rom_data[419]=rom_data[12];
    rom_data[420]=8'b01000100;
    rom_data[421]=rom_data[12];
    rom_data[422]=8'b01000100;
    rom_data[423]=rom_data[12];
    rom_data[424]=8'b01000100;
    rom_data[425]=rom_data[12];
    rom_data[426]=8'b01000100;
    rom_data[427]=rom_data[12];
    rom_data[428]=8'b01000100;
    rom_data[429]=rom_data[12];
    rom_data[430]=8'b01000101;
    rom_data[431]=rom_data[12];
    rom_data[432]=8'b01000101;
    rom_data[433]=rom_data[12];
    rom_data[434]=8'b01000101;
    rom_data[435]=rom_data[12];
    rom_data[436]=8'b01000101;
    rom_data[437]=rom_data[12];
    rom_data[438]=8'b01000101;
    rom_data[439]=rom_data[12];
    rom_data[440]=8'b01000101;
    rom_data[441]=rom_data[12];
    rom_data[442]=8'b01000101;
    rom_data[443]=rom_data[12];
    rom_data[444]=8'b01000110;
    rom_data[445]=rom_data[12];
    rom_data[446]=8'b01000110;
    rom_data[447]=rom_data[12];
    rom_data[448]=8'b01000110;
    rom_data[449]=rom_data[12];
    rom_data[450]=8'b01000110;
    rom_data[451]=rom_data[12];
    rom_data[452]=8'b01000110;
    rom_data[453]=rom_data[12];
    rom_data[454]=8'b01000110;
    rom_data[455]=rom_data[12];
    rom_data[456]=8'b01000110;
    rom_data[457]=rom_data[12];
    rom_data[458]=8'b01000111;
    rom_data[459]=rom_data[12];
    rom_data[460]=8'b01000111;
    rom_data[461]=rom_data[12];
    rom_data[462]=8'b01000111;
    rom_data[463]=rom_data[12];
    rom_data[464]=8'b01000111;
    rom_data[465]=rom_data[12];
    rom_data[466]=8'b01000111;
    rom_data[467]=rom_data[12];
    rom_data[468]=8'b01000111;
    rom_data[469]=rom_data[12];
    rom_data[470]=8'b01000111;
    rom_data[471]=rom_data[12];
    rom_data[472]=8'b01000111;
    rom_data[473]=rom_data[12];
    rom_data[474]=8'b01001000;
    rom_data[475]=rom_data[12];
    rom_data[476]=8'b01001000;
    rom_data[477]=rom_data[12];
    rom_data[478]=8'b01001000;
    rom_data[479]=rom_data[12];
    rom_data[480]=8'b01001000;
    rom_data[481]=rom_data[12];
    rom_data[482]=8'b01001000;
    rom_data[483]=rom_data[12];
    rom_data[484]=8'b01001000;
    rom_data[485]=rom_data[12];
    rom_data[486]=8'b01001000;
    rom_data[487]=rom_data[12];
    rom_data[488]=8'b01001000;
    rom_data[489]=rom_data[12];
    rom_data[490]=8'b01001001;
    rom_data[491]=rom_data[12];
    rom_data[492]=8'b01001001;
    rom_data[493]=rom_data[12];
    rom_data[494]=8'b01001001;
    rom_data[495]=rom_data[12];
    rom_data[496]=8'b01001001;
    rom_data[497]=rom_data[12];
    rom_data[498]=8'b01001001;
    rom_data[499]=rom_data[12];
    rom_data[500]=8'b01001001;
    rom_data[501]=rom_data[12];
    rom_data[502]=8'b01001001;
    rom_data[503]=rom_data[12];
    rom_data[504]=8'b01001001;
    rom_data[505]=rom_data[12];
    rom_data[506]=8'b01001001;
    rom_data[507]=rom_data[12];
    rom_data[508]=8'b01001010;
    rom_data[509]=rom_data[12];
    rom_data[510]=8'b01001010;
    rom_data[511]=rom_data[12];
    rom_data[512]=8'b01001010;
    rom_data[513]=rom_data[12];
    rom_data[514]=8'b01001010;
    rom_data[515]=rom_data[12];
    rom_data[516]=8'b01001010;
    rom_data[517]=rom_data[12];
    rom_data[518]=8'b01001010;
    rom_data[519]=rom_data[12];
    rom_data[520]=8'b01001010;
    rom_data[521]=rom_data[12];
    rom_data[522]=8'b01001010;
    rom_data[523]=rom_data[12];
    rom_data[524]=8'b01001010;
    rom_data[525]=rom_data[12];
    rom_data[526]=8'b01001011;
    rom_data[527]=rom_data[12];
    rom_data[528]=8'b01001011;
    rom_data[529]=rom_data[12];
    rom_data[530]=8'b01001011;
    rom_data[531]=rom_data[12];
    rom_data[532]=8'b01001011;
    rom_data[533]=rom_data[12];
    rom_data[534]=8'b01001011;
    rom_data[535]=rom_data[12];
    rom_data[536]=8'b01001011;
    rom_data[537]=rom_data[12];
    rom_data[538]=8'b01001011;
    rom_data[539]=rom_data[12];
    rom_data[540]=8'b01001011;
    rom_data[541]=rom_data[12];
    rom_data[542]=8'b01001011;
    rom_data[543]=rom_data[12];
    rom_data[544]=8'b01001011;
    rom_data[545]=rom_data[12];
    rom_data[546]=8'b01001100;
    rom_data[547]=rom_data[12];
    rom_data[548]=8'b01001100;
    rom_data[549]=rom_data[12];
    rom_data[550]=8'b01001100;
    rom_data[551]=rom_data[12];
    rom_data[552]=8'b01001100;
    rom_data[553]=rom_data[12];
    rom_data[554]=8'b01001100;
    rom_data[555]=rom_data[12];
    rom_data[556]=8'b01001100;
    rom_data[557]=rom_data[12];
    rom_data[558]=8'b01001100;
    rom_data[559]=rom_data[12];
    rom_data[560]=8'b01001100;
    rom_data[561]=rom_data[12];
    rom_data[562]=8'b01001100;
    rom_data[563]=rom_data[12];
    rom_data[564]=8'b01001100;
    rom_data[565]=rom_data[12];
    rom_data[566]=8'b01001101;
    rom_data[567]=rom_data[12];
    rom_data[568]=8'b01001101;
    rom_data[569]=rom_data[12];
    rom_data[570]=8'b01001101;
    rom_data[571]=rom_data[12];
    rom_data[572]=8'b01001101;
    rom_data[573]=rom_data[12];
    rom_data[574]=8'b01001101;
    rom_data[575]=rom_data[12];
    rom_data[576]=8'b01001101;
    rom_data[577]=rom_data[12];
    rom_data[578]=8'b01001101;
    rom_data[579]=rom_data[12];
    rom_data[580]=8'b01001101;
    rom_data[581]=rom_data[12];
    rom_data[582]=8'b01001101;
    rom_data[583]=rom_data[12];
    rom_data[584]=8'b01001101;
    rom_data[585]=rom_data[12];
    rom_data[586]=8'b01001110;
    rom_data[587]=rom_data[12];
    rom_data[588]=8'b01001110;
    rom_data[589]=rom_data[12];
    rom_data[590]=8'b01001110;
    rom_data[591]=rom_data[12];
    rom_data[592]=8'b01001110;
    rom_data[593]=rom_data[12];
    rom_data[594]=8'b01001110;
    rom_data[595]=rom_data[12];
    rom_data[596]=8'b01001110;
    rom_data[597]=rom_data[12];
    rom_data[598]=8'b01001110;
    rom_data[599]=rom_data[12];
    rom_data[600]=8'b01001110;
    rom_data[601]=rom_data[12];
    rom_data[602]=8'b01001111;
    rom_data[603]=rom_data[12];
    rom_data[604]=8'b01001111;
    rom_data[605]=rom_data[12];
    rom_data[606]=8'b01001111;
    rom_data[607]=rom_data[12];
    rom_data[608]=8'b01001111;
    rom_data[609]=rom_data[12];
    rom_data[610]=8'b01001111;
    rom_data[611]=rom_data[12];
    rom_data[612]=8'b01001111;
    rom_data[613]=rom_data[12];
    rom_data[614]=8'b01001111;
    rom_data[615]=rom_data[12];
    rom_data[616]=8'b01001111;
    rom_data[617]=rom_data[12];
    rom_data[618]=8'b01010000;
    rom_data[619]=rom_data[12];
    rom_data[620]=8'b01010000;
    rom_data[621]=rom_data[12];
    rom_data[622]=8'b01010000;
    rom_data[623]=rom_data[12];
    rom_data[624]=8'b01010000;
    rom_data[625]=rom_data[12];
    rom_data[626]=8'b01010000;
    rom_data[627]=rom_data[12];
    rom_data[628]=8'b01010000;
    rom_data[629]=rom_data[12];
    rom_data[630]=8'b01010000;
    rom_data[631]=rom_data[12];
    rom_data[632]=8'b01010001;
    rom_data[633]=rom_data[12];
    rom_data[634]=8'b01010001;
    rom_data[635]=rom_data[12];
    rom_data[636]=8'b01010001;
    rom_data[637]=rom_data[12];
    rom_data[638]=8'b01010001;
    rom_data[639]=rom_data[12];
    rom_data[640]=8'b01010001;
    rom_data[641]=rom_data[12];
    rom_data[642]=8'b01010001;
    rom_data[643]=rom_data[12];
    rom_data[644]=8'b01010001;
    rom_data[645]=rom_data[12];
    rom_data[646]=8'b01010001;
    rom_data[647]=rom_data[12];
    rom_data[648]=8'b01010010;
    rom_data[649]=rom_data[12];
    rom_data[650]=8'b01010010;
    rom_data[651]=rom_data[12];
    rom_data[652]=8'b01010010;
    rom_data[653]=rom_data[12];
    rom_data[654]=8'b01010010;
    rom_data[655]=rom_data[12];
    rom_data[656]=8'b01010010;
    rom_data[657]=rom_data[12];
    rom_data[658]=8'b01010010;
    rom_data[659]=rom_data[12];
    rom_data[660]=8'b01010010;
    rom_data[661]=rom_data[12];
    rom_data[662]=8'b01010011;
    rom_data[663]=rom_data[12];
    rom_data[664]=8'b01010011;
    rom_data[665]=rom_data[12];
    rom_data[666]=8'b01010011;
    rom_data[667]=rom_data[12];
    rom_data[668]=8'b01010011;
    rom_data[669]=rom_data[12];
    rom_data[670]=8'b01010011;
    rom_data[671]=rom_data[12];
    rom_data[672]=8'b01010011;
    rom_data[673]=rom_data[12];
    rom_data[674]=8'b01010011;
    rom_data[675]=rom_data[12];
    rom_data[676]=8'b01010011;
    rom_data[677]=rom_data[12];
    rom_data[678]=8'b01010011;
    rom_data[679]=rom_data[12];
    rom_data[680]=8'b01010100;
    rom_data[681]=rom_data[12];
    rom_data[682]=8'b01010100;
    rom_data[683]=rom_data[12];
    rom_data[684]=8'b01010100;
    rom_data[685]=rom_data[12];
    rom_data[686]=8'b01010100;
    rom_data[687]=rom_data[12];
    rom_data[688]=8'b01010100;
    rom_data[689]=rom_data[12];
    rom_data[690]=8'b01010100;
    rom_data[691]=rom_data[12];
    rom_data[692]=8'b01010100;
    rom_data[693]=rom_data[12];
    rom_data[694]=8'b01010100;
    rom_data[695]=rom_data[12];
    rom_data[696]=8'b01010100;
    rom_data[697]=rom_data[12];
    rom_data[698]=8'b01010101;
    rom_data[699]=rom_data[12];
    rom_data[700]=8'b01010101;
    rom_data[701]=rom_data[12];
    rom_data[702]=8'b01010101;
    rom_data[703]=rom_data[12];
    rom_data[704]=8'b01010101;
    rom_data[705]=rom_data[12];
    rom_data[706]=8'b01010101;
    rom_data[707]=rom_data[12];
    rom_data[708]=8'b01010101;
    rom_data[709]=rom_data[12];
    rom_data[710]=8'b01010101;
    rom_data[711]=rom_data[12];
    rom_data[712]=8'b01010101;
    rom_data[713]=rom_data[12];
    rom_data[714]=8'b01010101;
    rom_data[715]=rom_data[12];
    rom_data[716]=8'b01010101;
    rom_data[717]=rom_data[12];
    rom_data[718]=8'b01010110;
    rom_data[719]=rom_data[12];
    rom_data[720]=8'b01010110;
    rom_data[721]=rom_data[12];
    rom_data[722]=8'b01010110;
    rom_data[723]=rom_data[12];
    rom_data[724]=8'b01010110;
    rom_data[725]=rom_data[12];
    rom_data[726]=8'b01010110;
    rom_data[727]=rom_data[12];
    rom_data[728]=8'b01010110;
    rom_data[729]=rom_data[12];
    rom_data[730]=8'b01010110;
    rom_data[731]=rom_data[12];
    rom_data[732]=8'b01010110;
    rom_data[733]=rom_data[12];
    rom_data[734]=8'b01010110;
    rom_data[735]=rom_data[12];
    rom_data[736]=8'b01010110;
    rom_data[737]=rom_data[12];
    rom_data[738]=8'b01010111;
    rom_data[739]=rom_data[12];
    rom_data[740]=8'b01010111;
    rom_data[741]=rom_data[12];
    rom_data[742]=8'b01010111;
    rom_data[743]=rom_data[12];
    rom_data[744]=8'b01010111;
    rom_data[745]=rom_data[12];
    rom_data[746]=8'b01010111;
    rom_data[747]=rom_data[12];
    rom_data[748]=8'b01010111;
    rom_data[749]=rom_data[12];
    rom_data[750]=8'b01010111;
    rom_data[751]=rom_data[12];
    rom_data[752]=8'b01010111;
    rom_data[753]=rom_data[12];
    rom_data[754]=8'b01010111;
    rom_data[755]=rom_data[12];
    rom_data[756]=8'b01010111;
    rom_data[757]=rom_data[12];
    rom_data[758]=8'b01011000;
    rom_data[759]=rom_data[12];
    rom_data[760]=8'b01011000;
    rom_data[761]=rom_data[12];
    rom_data[762]=8'b01011000;
    rom_data[763]=rom_data[12];
    rom_data[764]=8'b01011000;
    rom_data[765]=rom_data[12];
    rom_data[766]=8'b01011000;
    rom_data[767]=rom_data[12];
    rom_data[768]=8'b01011000;
    rom_data[769]=rom_data[12];
    rom_data[770]=8'b01011000;
    rom_data[771]=rom_data[12];
    rom_data[772]=8'b01011000;
    rom_data[773]=rom_data[12];
    rom_data[774]=8'b01011000;
    rom_data[775]=rom_data[12];
    rom_data[776]=8'b01011001;
    rom_data[777]=rom_data[12];
    rom_data[778]=8'b01011001;
    rom_data[779]=rom_data[12];
    rom_data[780]=8'b01011001;
    rom_data[781]=rom_data[12];
    rom_data[782]=8'b01011001;
    rom_data[783]=rom_data[12];
    rom_data[784]=8'b01011001;
    rom_data[785]=rom_data[12];
    rom_data[786]=8'b01011001;
    rom_data[787]=rom_data[12];
    rom_data[788]=8'b01011001;
    rom_data[789]=rom_data[12];
    rom_data[790]=8'b01011001;
    rom_data[791]=rom_data[12];
    rom_data[792]=8'b01011010;
    rom_data[793]=rom_data[12];
    rom_data[794]=8'b01011010;
    rom_data[795]=rom_data[12];
    rom_data[796]=8'b01011010;
    rom_data[797]=rom_data[12];
    rom_data[798]=8'b01011010;
    rom_data[799]=rom_data[12];
    rom_data[800]=8'b01011010;
    rom_data[801]=rom_data[12];
    rom_data[802]=8'b01011010;
    rom_data[803]=rom_data[12];
    rom_data[804]=8'b01011010;
    rom_data[805]=rom_data[12];
    rom_data[806]=8'b01011011;
    rom_data[807]=rom_data[12];
    rom_data[808]=8'b01011011;
    rom_data[809]=rom_data[12];
    rom_data[810]=8'b01011011;
    rom_data[811]=rom_data[12];
    rom_data[812]=8'b01011011;
    rom_data[813]=rom_data[12];
    rom_data[814]=8'b01011011;
    rom_data[815]=rom_data[12];
    rom_data[816]=8'b01011011;
    rom_data[817]=rom_data[12];
    rom_data[818]=8'b01011011;
    rom_data[819]=rom_data[12];
    rom_data[820]=8'b01011011;
    rom_data[821]=rom_data[12];
    rom_data[822]=8'b01011100;
    rom_data[823]=rom_data[12];
    rom_data[824]=8'b01011100;
    rom_data[825]=rom_data[12];
    rom_data[826]=8'b01011100;
    rom_data[827]=rom_data[12];
    rom_data[828]=8'b01011100;
    rom_data[829]=rom_data[12];
    rom_data[830]=8'b01011100;
    rom_data[831]=rom_data[12];
    rom_data[832]=8'b01011100;
    rom_data[833]=rom_data[12];
    rom_data[834]=8'b01011100;
    rom_data[835]=rom_data[12];
    rom_data[836]=8'b01011101;
    rom_data[837]=rom_data[12];
    rom_data[838]=8'b01011101;
    rom_data[839]=rom_data[12];
    rom_data[840]=8'b01011101;
    rom_data[841]=rom_data[12];
    rom_data[842]=8'b01011101;
    rom_data[843]=rom_data[12];
    rom_data[844]=8'b01011101;
    rom_data[845]=rom_data[12];
    rom_data[846]=8'b01011101;
    rom_data[847]=rom_data[12];
    rom_data[848]=8'b01011101;
    rom_data[849]=rom_data[12];
    rom_data[850]=8'b01011101;
    rom_data[851]=rom_data[12];
    rom_data[852]=8'b01011110;
    rom_data[853]=rom_data[12];
    rom_data[854]=8'b01011110;
    rom_data[855]=rom_data[12];
    rom_data[856]=8'b01011110;
    rom_data[857]=rom_data[12];
    rom_data[858]=8'b01011110;
    rom_data[859]=rom_data[12];
    rom_data[860]=8'b01011110;
    rom_data[861]=rom_data[12];
    rom_data[862]=8'b01011110;
    rom_data[863]=rom_data[12];
    rom_data[864]=8'b01011110;
    rom_data[865]=rom_data[12];
    rom_data[866]=8'b01011110;
    rom_data[867]=rom_data[12];
    rom_data[868]=8'b01011110;
    rom_data[869]=rom_data[12];
    rom_data[870]=8'b01011111;
    rom_data[871]=rom_data[12];
    rom_data[872]=8'b01011111;
    rom_data[873]=rom_data[12];
    rom_data[874]=8'b01011111;
    rom_data[875]=rom_data[12];
    rom_data[876]=8'b01011111;
    rom_data[877]=rom_data[12];
    rom_data[878]=8'b01011111;
    rom_data[879]=rom_data[12];
    rom_data[880]=8'b01011111;
    rom_data[881]=rom_data[12];
    rom_data[882]=8'b01011111;
    rom_data[883]=rom_data[12];
    rom_data[884]=8'b01011111;
    rom_data[885]=rom_data[12];
    rom_data[886]=8'b01011111;
    rom_data[887]=rom_data[12];
    rom_data[888]=8'b01011111;
    rom_data[889]=rom_data[12];
    rom_data[890]=8'b01100000;
    rom_data[891]=rom_data[12];
    rom_data[892]=8'b01100000;
    rom_data[893]=rom_data[12];
    rom_data[894]=8'b01100000;
    rom_data[895]=rom_data[12];
    rom_data[896]=8'b01100000;
    rom_data[897]=rom_data[12];
    rom_data[898]=8'b01100000;
    rom_data[899]=rom_data[12];
    rom_data[900]=8'b01100000;
    rom_data[901]=rom_data[12];
    rom_data[902]=8'b01100000;
    rom_data[903]=rom_data[12];
    rom_data[904]=8'b01100000;
    rom_data[905]=rom_data[12];
    rom_data[906]=8'b01100000;
    rom_data[907]=rom_data[12];
    rom_data[908]=8'b01100000;
    rom_data[909]=rom_data[12];
    rom_data[910]=8'b01100001;
    rom_data[911]=rom_data[12];
    rom_data[912]=8'b01100001;
    rom_data[913]=rom_data[12];
    rom_data[914]=8'b01100001;
    rom_data[915]=rom_data[12];
    rom_data[916]=8'b01100001;
    rom_data[917]=rom_data[12];
    rom_data[918]=8'b01100001;
    rom_data[919]=rom_data[12];
    rom_data[920]=8'b01100001;
    rom_data[921]=rom_data[12];
    rom_data[922]=8'b01100001;
    rom_data[923]=rom_data[12];
    rom_data[924]=8'b01100001;
    rom_data[925]=rom_data[12];
    rom_data[926]=8'b01100001;
    rom_data[927]=rom_data[12];
    rom_data[928]=8'b01100001;
    rom_data[929]=rom_data[12];
    rom_data[930]=8'b01100010;
    rom_data[931]=rom_data[12];
    rom_data[932]=8'b01100010;
    rom_data[933]=rom_data[12];
    rom_data[934]=8'b01100010;
    rom_data[935]=rom_data[12];
    rom_data[936]=8'b01100010;
    rom_data[937]=rom_data[12];
    rom_data[938]=8'b01100010;
    rom_data[939]=rom_data[12];
    rom_data[940]=8'b01100010;
    rom_data[941]=rom_data[12];
    rom_data[942]=8'b01100010;
    rom_data[943]=rom_data[12];
    rom_data[944]=8'b01100010;
    rom_data[945]=rom_data[12];
    rom_data[946]=8'b01100010;
    rom_data[947]=rom_data[12];
    rom_data[948]=8'b01100011;
    rom_data[949]=rom_data[12];
    rom_data[950]=8'b01100011;
    rom_data[951]=rom_data[12];
    rom_data[952]=8'b01100011;
    rom_data[953]=rom_data[12];
    rom_data[954]=8'b01100011;
    rom_data[955]=rom_data[12];
    rom_data[956]=8'b01100011;
    rom_data[957]=rom_data[12];
    rom_data[958]=8'b01100011;
    rom_data[959]=rom_data[12];
    rom_data[960]=8'b01100011;
    rom_data[961]=rom_data[12];
    rom_data[962]=8'b01100011;
    rom_data[963]=rom_data[12];
    rom_data[964]=8'b01100011;
    rom_data[965]=rom_data[12];
    rom_data[966]=8'b01100100;
    rom_data[967]=rom_data[12];
    rom_data[968]=8'b01100100;
    rom_data[969]=rom_data[12];
    rom_data[970]=8'b01100100;
    rom_data[971]=rom_data[12];
    rom_data[972]=8'b01100100;
    rom_data[973]=rom_data[12];
    rom_data[974]=8'b01100100;
    rom_data[975]=rom_data[12];
    rom_data[976]=8'b01100100;
    rom_data[977]=rom_data[12];
    rom_data[978]=8'b01100100;
    rom_data[979]=rom_data[12];
    rom_data[980]=8'b01100101;
    rom_data[981]=rom_data[12];
    rom_data[982]=8'b01100101;
    rom_data[983]=rom_data[12];
    rom_data[984]=8'b01100101;
    rom_data[985]=rom_data[12];
    rom_data[986]=8'b01100101;
    rom_data[987]=rom_data[12];
    rom_data[988]=8'b01100101;
    rom_data[989]=rom_data[12];
    rom_data[990]=8'b01100101;
    rom_data[991]=rom_data[12];
    rom_data[992]=8'b01100101;
    rom_data[993]=rom_data[12];
    rom_data[994]=8'b01100110;
    rom_data[995]=rom_data[12];
    rom_data[996]=8'b01100110;
    rom_data[997]=rom_data[12];
    rom_data[998]=8'b01100110;
    rom_data[999]=rom_data[12];
    rom_data[1000]=8'b01100110;
    rom_data[1001]=rom_data[12];
    rom_data[1002]=8'b01100110;
    rom_data[1003]=rom_data[12];
    rom_data[1004]=8'b01100110;
    rom_data[1005]=rom_data[12];
    rom_data[1006]=8'b01100110;
    rom_data[1007]=rom_data[12];
    rom_data[1008]=8'b01100110;
    rom_data[1009]=rom_data[12];
    rom_data[1010]=8'b01100111;
    rom_data[1011]=rom_data[12];
    rom_data[1012]=8'b01100111;
    rom_data[1013]=rom_data[12];
    rom_data[1014]=8'b01100111;
    rom_data[1015]=rom_data[12];
    rom_data[1016]=8'b01100111;
    rom_data[1017]=rom_data[12];
    rom_data[1018]=8'b01100111;
    rom_data[1019]=rom_data[12];
    rom_data[1020]=8'b01100111;
    rom_data[1021]=rom_data[12];
    rom_data[1022]=8'b01100111;
    rom_data[1023]=rom_data[12];
    rom_data[1024]=8'b01101000;
    rom_data[1025]=rom_data[12];
    rom_data[1026]=8'b01101000;
    rom_data[1027]=rom_data[12];
    rom_data[1028]=8'b01101000;
    rom_data[1029]=rom_data[12];
    rom_data[1030]=8'b01101000;
    rom_data[1031]=rom_data[12];
    rom_data[1032]=8'b01101000;
    rom_data[1033]=rom_data[12];
    rom_data[1034]=8'b01101000;
    rom_data[1035]=rom_data[12];
    rom_data[1036]=8'b01101000;
    rom_data[1037]=rom_data[12];
    rom_data[1038]=8'b01101000;
    rom_data[1039]=rom_data[12];
    rom_data[1040]=8'b01101000;
    rom_data[1041]=rom_data[12];
    rom_data[1042]=8'b01101001;
    rom_data[1043]=rom_data[12];
    rom_data[1044]=8'b01101001;
    rom_data[1045]=rom_data[12];
    rom_data[1046]=8'b01101001;
    rom_data[1047]=rom_data[12];
    rom_data[1048]=8'b01101001;
    rom_data[1049]=rom_data[12];
    rom_data[1050]=8'b01101001;
    rom_data[1051]=rom_data[12];
    rom_data[1052]=8'b01101001;
    rom_data[1053]=rom_data[12];
    rom_data[1054]=8'b01101001;
    rom_data[1055]=rom_data[12];
    rom_data[1056]=8'b01101001;
    rom_data[1057]=rom_data[12];
    rom_data[1058]=8'b01101001;
    rom_data[1059]=rom_data[12];
    rom_data[1060]=8'b01101001;
    rom_data[1061]=rom_data[12];
    rom_data[1062]=8'b01101010;
    rom_data[1063]=rom_data[12];
    rom_data[1064]=8'b01101010;
    rom_data[1065]=rom_data[12];
    rom_data[1066]=8'b01101010;
    rom_data[1067]=rom_data[12];
    rom_data[1068]=8'b01101010;
    rom_data[1069]=rom_data[12];
    rom_data[1070]=8'b01101010;
    rom_data[1071]=rom_data[12];
    rom_data[1072]=8'b01101010;
    rom_data[1073]=rom_data[12];
    rom_data[1074]=8'b01101010;
    rom_data[1075]=rom_data[12];
    rom_data[1076]=8'b01101010;
    rom_data[1077]=rom_data[12];
    rom_data[1078]=8'b01101010;
    rom_data[1079]=rom_data[12];
    rom_data[1080]=8'b01101011;
    rom_data[1081]=rom_data[12];
    rom_data[1082]=8'b01101011;
    rom_data[1083]=rom_data[12];
    rom_data[1084]=8'b01101011;
    rom_data[1085]=rom_data[12];
    rom_data[1086]=8'b01101011;
    rom_data[1087]=rom_data[12];
    rom_data[1088]=8'b01101011;
    rom_data[1089]=rom_data[12];
    rom_data[1090]=8'b01101011;
    rom_data[1091]=rom_data[12];
    rom_data[1092]=8'b01101011;
    rom_data[1093]=rom_data[12];
    rom_data[1094]=8'b01101011;
    rom_data[1095]=rom_data[12];
    rom_data[1096]=8'b01101011;
    rom_data[1097]=rom_data[12];
    rom_data[1098]=8'b01101011;
    rom_data[1099]=rom_data[12];
    rom_data[1100]=8'b01101100;
    rom_data[1101]=rom_data[12];
    rom_data[1102]=8'b01101100;
    rom_data[1103]=rom_data[12];
    rom_data[1104]=8'b01101100;
    rom_data[1105]=rom_data[12];
    rom_data[1106]=8'b01101100;
    rom_data[1107]=rom_data[12];
    rom_data[1108]=8'b01101100;
    rom_data[1109]=rom_data[12];
    rom_data[1110]=8'b01101100;
    rom_data[1111]=rom_data[12];
    rom_data[1112]=8'b01101100;
    rom_data[1113]=rom_data[12];
    rom_data[1114]=8'b01101100;
    rom_data[1115]=rom_data[12];
    rom_data[1116]=8'b01101100;
    rom_data[1117]=rom_data[12];
    rom_data[1118]=8'b01101100;
    rom_data[1119]=rom_data[12];
    rom_data[1120]=8'b01101101;
    rom_data[1121]=rom_data[12];
    rom_data[1122]=8'b01101101;
    rom_data[1123]=rom_data[12];
    rom_data[1124]=8'b01101101;
    rom_data[1125]=rom_data[12];
    rom_data[1126]=8'b01101101;
    rom_data[1127]=rom_data[12];
    rom_data[1128]=8'b01101101;
    rom_data[1129]=rom_data[12];
    rom_data[1130]=8'b01101101;
    rom_data[1131]=rom_data[12];
    rom_data[1132]=8'b01101101;
    rom_data[1133]=rom_data[12];
    rom_data[1134]=8'b01101101;
    rom_data[1135]=rom_data[12];
    rom_data[1136]=8'b01101101;
    rom_data[1137]=rom_data[12];
    rom_data[1138]=8'b01101110;
    rom_data[1139]=rom_data[12];
    rom_data[1140]=8'b01101110;
    rom_data[1141]=rom_data[12];
    rom_data[1142]=8'b01101110;
    rom_data[1143]=rom_data[12];
    rom_data[1144]=8'b01101110;
    rom_data[1145]=rom_data[12];
    rom_data[1146]=8'b01101110;
    rom_data[1147]=rom_data[12];
    rom_data[1148]=8'b01101110;
    rom_data[1149]=rom_data[12];
    rom_data[1150]=8'b01101110;
    rom_data[1151]=rom_data[12];
    rom_data[1152]=8'b01101110;
    rom_data[1153]=rom_data[12];
    rom_data[1154]=8'b01101111;
    rom_data[1155]=rom_data[12];
    rom_data[1156]=8'b01101111;
    rom_data[1157]=rom_data[12];
    rom_data[1158]=8'b01101111;
    rom_data[1159]=rom_data[12];
    rom_data[1160]=8'b01101111;
    rom_data[1161]=rom_data[12];
    rom_data[1162]=8'b01101111;
    rom_data[1163]=rom_data[12];
    rom_data[1164]=8'b01101111;
    rom_data[1165]=rom_data[12];
    rom_data[1166]=8'b01101111;
    rom_data[1167]=rom_data[12];
    rom_data[1168]=8'b01110000;
    rom_data[1169]=rom_data[12];
    rom_data[1170]=8'b01110000;
    rom_data[1171]=rom_data[12];
    rom_data[1172]=8'b01110000;
    rom_data[1173]=rom_data[12];
    rom_data[1174]=8'b01110000;
    rom_data[1175]=rom_data[12];
    rom_data[1176]=8'b01110000;
    rom_data[1177]=rom_data[12];
    rom_data[1178]=8'b01110000;
    rom_data[1179]=rom_data[12];
    rom_data[1180]=8'b01110000;
    rom_data[1181]=rom_data[12];
    rom_data[1182]=8'b01110000;
    rom_data[1183]=rom_data[12];
    rom_data[1184]=8'b01110001;
    rom_data[1185]=rom_data[12];
    rom_data[1186]=8'b01110001;
    rom_data[1187]=rom_data[12];
    rom_data[1188]=8'b01110001;
    rom_data[1189]=rom_data[12];
    rom_data[1190]=8'b01110001;
    rom_data[1191]=rom_data[12];
    rom_data[1192]=8'b01110001;
    rom_data[1193]=rom_data[12];
    rom_data[1194]=8'b01110001;
    rom_data[1195]=rom_data[12];
    rom_data[1196]=8'b01110001;
    rom_data[1197]=rom_data[12];
    rom_data[1198]=8'b01110010;
    rom_data[1199]=rom_data[12];
    rom_data[1200]=8'b01110010;
    rom_data[1201]=rom_data[12];
    rom_data[1202]=8'b01110010;
    rom_data[1203]=rom_data[12];
    rom_data[1204]=8'b01110010;
    rom_data[1205]=rom_data[12];
    rom_data[1206]=8'b01110010;
    rom_data[1207]=rom_data[12];
    rom_data[1208]=8'b01110010;
    rom_data[1209]=rom_data[12];
    rom_data[1210]=8'b01110010;
    rom_data[1211]=rom_data[12];
    rom_data[1212]=8'b01110010;
    rom_data[1213]=rom_data[12];
    rom_data[1214]=8'b01110011;
    rom_data[1215]=rom_data[12];
    rom_data[1216]=8'b01110011;
    rom_data[1217]=rom_data[12];
    rom_data[1218]=8'b01110011;
    rom_data[1219]=rom_data[12];
    rom_data[1220]=8'b01110011;
    rom_data[1221]=rom_data[12];
    rom_data[1222]=8'b01110011;
    rom_data[1223]=rom_data[12];
    rom_data[1224]=8'b01110011;
    rom_data[1225]=rom_data[12];
    rom_data[1226]=8'b01110011;
    rom_data[1227]=rom_data[12];
    rom_data[1228]=8'b01110011;
    rom_data[1229]=rom_data[12];
    rom_data[1230]=8'b01110011;
    rom_data[1231]=rom_data[12];
    rom_data[1232]=8'b01110100;
    rom_data[1233]=rom_data[12];
    rom_data[1234]=8'b01110100;
    rom_data[1235]=rom_data[12];
    rom_data[1236]=8'b01110100;
    rom_data[1237]=rom_data[12];
    rom_data[1238]=8'b01110100;
    rom_data[1239]=rom_data[12];
    rom_data[1240]=8'b01110100;
    rom_data[1241]=rom_data[12];
    rom_data[1242]=8'b01110100;
    rom_data[1243]=rom_data[12];
    rom_data[1244]=8'b01110100;
    rom_data[1245]=rom_data[12];
    rom_data[1246]=8'b01110100;
    rom_data[1247]=rom_data[12];
    rom_data[1248]=8'b01110100;
    rom_data[1249]=rom_data[12];
    rom_data[1250]=8'b01110100;
    rom_data[1251]=rom_data[12];
    rom_data[1252]=8'b01110101;
    rom_data[1253]=rom_data[12];
    rom_data[1254]=8'b01110101;
    rom_data[1255]=rom_data[12];
    rom_data[1256]=8'b01110101;
    rom_data[1257]=rom_data[12];
    rom_data[1258]=8'b01110101;
    rom_data[1259]=rom_data[12];
    rom_data[1260]=8'b01110101;
    rom_data[1261]=rom_data[12];
    rom_data[1262]=8'b01110101;
    rom_data[1263]=rom_data[12];
    rom_data[1264]=8'b01110101;
    rom_data[1265]=rom_data[12];
    rom_data[1266]=8'b01110101;
    rom_data[1267]=rom_data[12];
    rom_data[1268]=8'b01110101;
    rom_data[1269]=rom_data[12];
    rom_data[1270]=8'b01110101;
    rom_data[1271]=rom_data[12];
    rom_data[1272]=8'b01110110;
    rom_data[1273]=rom_data[12];
    rom_data[1274]=8'b01110110;
    rom_data[1275]=rom_data[12];
    rom_data[1276]=8'b01110110;
    rom_data[1277]=rom_data[12];
    rom_data[1278]=8'b01110110;
    rom_data[1279]=rom_data[12];
    rom_data[1280]=8'b01110110;
    rom_data[1281]=rom_data[12];
    rom_data[1282]=8'b01110110;
    rom_data[1283]=rom_data[12];
    rom_data[1284]=8'b01110110;
    rom_data[1285]=rom_data[12];
    rom_data[1286]=8'b01110110;
    rom_data[1287]=rom_data[12];
    rom_data[1288]=8'b01110110;
    rom_data[1289]=rom_data[12];
    rom_data[1290]=8'b01110110;
    rom_data[1291]=rom_data[12];
    rom_data[1292]=8'b01110111;
    rom_data[1293]=rom_data[12];
    rom_data[1294]=8'b01110111;
    rom_data[1295]=rom_data[12];
    rom_data[1296]=8'b01110111;
    rom_data[1297]=rom_data[12];
    rom_data[1298]=8'b01110111;
    rom_data[1299]=rom_data[12];
    rom_data[1300]=8'b01110111;
    rom_data[1301]=rom_data[12];
    rom_data[1302]=8'b01110111;
    rom_data[1303]=rom_data[12];
    rom_data[1304]=8'b01110111;
    rom_data[1305]=rom_data[12];
    rom_data[1306]=8'b01110111;
    rom_data[1307]=rom_data[12];
    rom_data[1308]=8'b01110111;
    rom_data[1309]=rom_data[12];
    rom_data[1310]=8'b01111000;
    rom_data[1311]=rom_data[12];
    rom_data[1312]=8'b01111000;
    rom_data[1313]=rom_data[12];
    rom_data[1314]=8'b01111000;
    rom_data[1315]=rom_data[12];
    rom_data[1316]=8'b01111000;
    rom_data[1317]=rom_data[12];
    rom_data[1318]=8'b01111000;
    rom_data[1319]=rom_data[12];
    rom_data[1320]=8'b01111000;
    rom_data[1321]=rom_data[12];
    rom_data[1322]=8'b01111000;
    rom_data[1323]=rom_data[12];
    rom_data[1324]=8'b01111000;
    rom_data[1325]=rom_data[12];
    rom_data[1326]=8'b01111000;
    rom_data[1327]=rom_data[12];
    rom_data[1328]=8'b01111001;
    rom_data[1329]=rom_data[12];
    rom_data[1330]=8'b01111001;
    rom_data[1331]=rom_data[12];
    rom_data[1332]=8'b01111001;
    rom_data[1333]=rom_data[12];
    rom_data[1334]=8'b01111001;
    rom_data[1335]=rom_data[12];
    rom_data[1336]=8'b01111001;
    rom_data[1337]=rom_data[12];
    rom_data[1338]=8'b01111001;
    rom_data[1339]=rom_data[12];
    rom_data[1340]=8'b01111001;
    rom_data[1341]=rom_data[12];
    rom_data[1342]=8'b01111010;
    rom_data[1343]=rom_data[12];
    rom_data[1344]=8'b01111010;
    rom_data[1345]=rom_data[12];
    rom_data[1346]=8'b01111010;
    rom_data[1347]=rom_data[12];
    rom_data[1348]=8'b01111010;
    rom_data[1349]=rom_data[12];
    rom_data[1350]=8'b01111010;
    rom_data[1351]=rom_data[12];
    rom_data[1352]=8'b01111010;
    rom_data[1353]=rom_data[12];
    rom_data[1354]=8'b01111010;
    rom_data[1355]=rom_data[12];
    rom_data[1356]=8'b01111011;
    rom_data[1357]=rom_data[12];
    rom_data[1358]=8'b01111011;
    rom_data[1359]=rom_data[12];
    rom_data[1360]=8'b01111011;
    rom_data[1361]=rom_data[12];
    rom_data[1362]=8'b01111011;
    rom_data[1363]=rom_data[12];
    rom_data[1364]=8'b01111011;
    rom_data[1365]=rom_data[12];
    rom_data[1366]=8'b01111011;
    rom_data[1367]=rom_data[12];
    rom_data[1368]=8'b01111011;
    rom_data[1369]=rom_data[12];
    rom_data[1370]=8'b01111011;
    rom_data[1371]=rom_data[12];
    rom_data[1372]=8'b01111100;
    rom_data[1373]=rom_data[12];
    rom_data[1374]=8'b01111100;
    rom_data[1375]=rom_data[12];
    rom_data[1376]=8'b01111100;
    rom_data[1377]=rom_data[12];
    rom_data[1378]=8'b01111100;
    rom_data[1379]=rom_data[12];
    rom_data[1380]=8'b01111100;
    rom_data[1381]=rom_data[12];
    rom_data[1382]=8'b01111100;
    rom_data[1383]=rom_data[12];
    rom_data[1384]=8'b01111100;
    rom_data[1385]=rom_data[12];
    rom_data[1386]=8'b01111100;
    rom_data[1387]=rom_data[12];
    rom_data[1388]=8'b01111101;
    rom_data[1389]=rom_data[12];
    rom_data[1390]=8'b01111101;
    rom_data[1391]=rom_data[12];
    rom_data[1392]=8'b01111101;
    rom_data[1393]=rom_data[12];
    rom_data[1394]=8'b01111101;
    rom_data[1395]=rom_data[12];
    rom_data[1396]=8'b01111101;
    rom_data[1397]=rom_data[12];
    rom_data[1398]=8'b01111101;
    rom_data[1399]=rom_data[12];
    rom_data[1400]=8'b01111101;
    rom_data[1401]=rom_data[12];
    rom_data[1402]=8'b01111101;
    rom_data[1403]=rom_data[12];
    rom_data[1404]=8'b01111110;
    rom_data[1405]=rom_data[12];
    rom_data[1406]=8'b01111110;
    rom_data[1407]=rom_data[12];
    rom_data[1408]=8'b01111110;
    rom_data[1409]=rom_data[12];
    rom_data[1410]=8'b01111110;
    rom_data[1411]=rom_data[12];
    rom_data[1412]=8'b01111110;
    rom_data[1413]=rom_data[12];
    rom_data[1414]=8'b01111110;
    rom_data[1415]=rom_data[12];
    rom_data[1416]=8'b01111110;
    rom_data[1417]=rom_data[12];
    rom_data[1418]=8'b01111110;
    rom_data[1419]=rom_data[12];
    rom_data[1420]=8'b01111110;
    rom_data[1421]=rom_data[12];
    rom_data[1422]=8'b01111110;
    rom_data[1423]=rom_data[12];
    rom_data[1424]=8'b01111111;
    rom_data[1425]=rom_data[12];
    rom_data[1426]=8'b01111111;
    rom_data[1427]=rom_data[12];
    rom_data[1428]=8'b01111111;
    rom_data[1429]=rom_data[12];
    rom_data[1430]=8'b01111111;
    rom_data[1431]=rom_data[12];
    rom_data[1432]=8'b01111111;
    rom_data[1433]=rom_data[12];
    rom_data[1434]=8'b01111111;
    rom_data[1435]=rom_data[12];
    rom_data[1436]=8'b01111111;
    rom_data[1437]=rom_data[12];
    rom_data[1438]=8'b01111111;
    rom_data[1439]=rom_data[12];
    rom_data[1440]=8'b01111111;
    rom_data[1441]=rom_data[12];
    rom_data[1442]=8'b01111111;
    rom_data[1443]=rom_data[12];
    rom_data[1444]=8'b10000000;
    rom_data[1445]=rom_data[12];
    rom_data[1446]=8'b10000000;
    rom_data[1447]=rom_data[12];
    rom_data[1448]=8'b10000000;
    rom_data[1449]=rom_data[12];
    rom_data[1450]=8'b10000000;
    rom_data[1451]=rom_data[12];
    rom_data[1452]=8'b10000000;
    rom_data[1453]=rom_data[12];
    rom_data[1454]=8'b10000000;
    rom_data[1455]=rom_data[12];
    rom_data[1456]=8'b10000000;
    rom_data[1457]=rom_data[12];
    rom_data[1458]=8'b10000000;
    rom_data[1459]=rom_data[12];
    rom_data[1460]=8'b10000000;
    rom_data[1461]=rom_data[12];
    rom_data[1462]=8'b10000000;
    rom_data[1463]=rom_data[12];
    rom_data[1464]=8'b10000001;
    rom_data[1465]=rom_data[12];
    rom_data[1466]=8'b10000001;
    rom_data[1467]=rom_data[12];
    rom_data[1468]=8'b10000001;
    rom_data[1469]=rom_data[12];
    rom_data[1470]=8'b10000001;
    rom_data[1471]=rom_data[12];
    rom_data[1472]=8'b10000001;
    rom_data[1473]=rom_data[12];
    rom_data[1474]=8'b10000001;
    rom_data[1475]=rom_data[12];
    rom_data[1476]=8'b10000001;
    rom_data[1477]=rom_data[12];
    rom_data[1478]=8'b10000001;
    rom_data[1479]=rom_data[12];
    rom_data[1480]=8'b10000001;
    rom_data[1481]=rom_data[12];
    rom_data[1482]=8'b10000010;
    rom_data[1483]=rom_data[12];
    rom_data[1484]=8'b10000010;
    rom_data[1485]=rom_data[12];
    rom_data[1486]=8'b10000010;
    rom_data[1487]=rom_data[12];
    rom_data[1488]=8'b10000010;
    rom_data[1489]=rom_data[12];
    rom_data[1490]=8'b10000010;
    rom_data[1491]=rom_data[12];
    rom_data[1492]=8'b10000010;
    rom_data[1493]=rom_data[12];
    rom_data[1494]=8'b10000010;
    rom_data[1495]=rom_data[12];
    rom_data[1496]=8'b10000010;
    rom_data[1497]=rom_data[12];
    rom_data[1498]=8'b10000010;
    rom_data[1499]=rom_data[12];
    rom_data[1500]=8'b10000011;
    rom_data[1501]=rom_data[12];
    rom_data[1502]=8'b10000011;
    rom_data[1503]=rom_data[12];
    rom_data[1504]=8'b10000011;
    rom_data[1505]=rom_data[12];
    rom_data[1506]=8'b10000011;
    rom_data[1507]=rom_data[12];
    rom_data[1508]=8'b10000011;
    rom_data[1509]=rom_data[12];
    rom_data[1510]=8'b10000011;
    rom_data[1511]=rom_data[12];
    rom_data[1512]=8'b10000011;
    rom_data[1513]=rom_data[12];
    rom_data[1514]=8'b10000011;
    rom_data[1515]=rom_data[12];
    rom_data[1516]=8'b10000100;
    rom_data[1517]=rom_data[12];
    rom_data[1518]=8'b10000100;
    rom_data[1519]=rom_data[12];
    rom_data[1520]=8'b10000100;
    rom_data[1521]=rom_data[12];
    rom_data[1522]=8'b10000100;
    rom_data[1523]=rom_data[12];
    rom_data[1524]=8'b10000100;
    rom_data[1525]=rom_data[12];
    rom_data[1526]=8'b10000100;
    rom_data[1527]=rom_data[12];
    rom_data[1528]=8'b10000100;
    rom_data[1529]=rom_data[12];
    rom_data[1530]=8'b10000101;
    rom_data[1531]=rom_data[12];
    rom_data[1532]=8'b10000101;
    rom_data[1533]=rom_data[12];
    rom_data[1534]=8'b10000101;
    rom_data[1535]=rom_data[12];
    rom_data[1536]=8'b10000101;
    rom_data[1537]=rom_data[12];
    rom_data[1538]=8'b10000101;
    rom_data[1539]=rom_data[12];
    rom_data[1540]=8'b10000101;
    rom_data[1541]=rom_data[12];
    rom_data[1542]=8'b10000101;
    rom_data[1543]=rom_data[12];
    rom_data[1544]=8'b10000101;
    rom_data[1545]=rom_data[12];
    rom_data[1546]=8'b10000110;
    rom_data[1547]=rom_data[12];
    rom_data[1548]=8'b10000110;
    rom_data[1549]=rom_data[12];
    rom_data[1550]=8'b10000110;
    rom_data[1551]=rom_data[12];
    rom_data[1552]=8'b10000110;
    rom_data[1553]=rom_data[12];
    rom_data[1554]=8'b10000110;
    rom_data[1555]=rom_data[12];
    rom_data[1556]=8'b10000110;
    rom_data[1557]=rom_data[12];
    rom_data[1558]=8'b10000110;
    rom_data[1559]=rom_data[12];
    rom_data[1560]=8'b10000111;
    rom_data[1561]=rom_data[12];
    rom_data[1562]=8'b10000111;
    rom_data[1563]=rom_data[12];
    rom_data[1564]=8'b10000111;
    rom_data[1565]=rom_data[12];
    rom_data[1566]=8'b10000111;
    rom_data[1567]=rom_data[12];
    rom_data[1568]=8'b10000111;
    rom_data[1569]=rom_data[12];
    rom_data[1570]=8'b10000111;
    rom_data[1571]=rom_data[12];
    rom_data[1572]=8'b10000111;
    rom_data[1573]=rom_data[12];
    rom_data[1574]=8'b10000111;
    rom_data[1575]=rom_data[12];
    rom_data[1576]=8'b10000111;
    rom_data[1577]=rom_data[12];
    rom_data[1578]=8'b10001000;
    rom_data[1579]=rom_data[12];
    rom_data[1580]=8'b10001000;
    rom_data[1581]=rom_data[12];
    rom_data[1582]=8'b10001000;
    rom_data[1583]=rom_data[12];
    rom_data[1584]=8'b10001000;
    rom_data[1585]=rom_data[12];
    rom_data[1586]=8'b10001000;
    rom_data[1587]=rom_data[12];
    rom_data[1588]=8'b10001000;
    rom_data[1589]=rom_data[12];
    rom_data[1590]=8'b10001000;
    rom_data[1591]=rom_data[12];
    rom_data[1592]=8'b10001000;
    rom_data[1593]=rom_data[12];
    rom_data[1594]=8'b10001000;
    rom_data[1595]=rom_data[12];
    rom_data[1596]=8'b10001001;
    rom_data[1597]=rom_data[12];
    rom_data[1598]=8'b10001001;
    rom_data[1599]=rom_data[12];
    rom_data[1600]=8'b10001001;
    rom_data[1601]=rom_data[12];
    rom_data[1602]=8'b10001001;
    rom_data[1603]=rom_data[12];
    rom_data[1604]=8'b10001001;
    rom_data[1605]=rom_data[12];
    rom_data[1606]=8'b10001001;
    rom_data[1607]=rom_data[12];
    rom_data[1608]=8'b10001001;
    rom_data[1609]=rom_data[12];
    rom_data[1610]=8'b10001001;
    rom_data[1611]=rom_data[12];
    rom_data[1612]=8'b10001001;
    rom_data[1613]=rom_data[12];
    rom_data[1614]=8'b10001001;
    rom_data[1615]=rom_data[12];
    rom_data[1616]=8'b10001010;
    rom_data[1617]=rom_data[12];
    rom_data[1618]=8'b10001010;
    rom_data[1619]=rom_data[12];
    rom_data[1620]=8'b10001010;
    rom_data[1621]=rom_data[12];
    rom_data[1622]=8'b10001010;
    rom_data[1623]=rom_data[12];
    rom_data[1624]=8'b10001010;
    rom_data[1625]=rom_data[12];
    rom_data[1626]=8'b10001010;
    rom_data[1627]=rom_data[12];
    rom_data[1628]=8'b10001001;
    rom_data[1629]=rom_data[12];
    rom_data[1630]=8'b10001001;
    rom_data[1631]=rom_data[12];
    rom_data[1632]=8'b10001001;
    rom_data[1633]=rom_data[12];
    rom_data[1634]=8'b10001001;
    rom_data[1635]=rom_data[12];
    rom_data[1636]=8'b10001001;
    rom_data[1637]=rom_data[12];
    rom_data[1638]=8'b10001001;
    rom_data[1639]=rom_data[12];
    rom_data[1640]=8'b10001001;
    rom_data[1641]=rom_data[12];
    rom_data[1642]=8'b10001001;
    rom_data[1643]=rom_data[12];
    rom_data[1644]=8'b10001001;
    rom_data[1645]=rom_data[12];
    rom_data[1646]=8'b10001001;
    rom_data[1647]=rom_data[12];
    rom_data[1648]=8'b10001000;
    rom_data[1649]=rom_data[12];
    rom_data[1650]=8'b10001000;
    rom_data[1651]=rom_data[12];
    rom_data[1652]=8'b10001000;
    rom_data[1653]=rom_data[12];
    rom_data[1654]=8'b10001000;
    rom_data[1655]=rom_data[12];
    rom_data[1656]=8'b10001000;
    rom_data[1657]=rom_data[12];
    rom_data[1658]=8'b10001000;
    rom_data[1659]=rom_data[12];
    rom_data[1660]=8'b10001000;
    rom_data[1661]=rom_data[12];
    rom_data[1662]=8'b10001000;
    rom_data[1663]=rom_data[12];
    rom_data[1664]=8'b10001000;
    rom_data[1665]=rom_data[12];
    rom_data[1666]=8'b10000111;
    rom_data[1667]=rom_data[12];
    rom_data[1668]=8'b10000111;
    rom_data[1669]=rom_data[12];
    rom_data[1670]=8'b10000111;
    rom_data[1671]=rom_data[12];
    rom_data[1672]=8'b10000111;
    rom_data[1673]=rom_data[12];
    rom_data[1674]=8'b10000111;
    rom_data[1675]=rom_data[12];
    rom_data[1676]=8'b10000111;
    rom_data[1677]=rom_data[12];
    rom_data[1678]=8'b10000111;
    rom_data[1679]=rom_data[12];
    rom_data[1680]=8'b10000111;
    rom_data[1681]=rom_data[12];
    rom_data[1682]=8'b10000111;
    rom_data[1683]=rom_data[12];
    rom_data[1684]=8'b10000110;
    rom_data[1685]=rom_data[12];
    rom_data[1686]=8'b10000110;
    rom_data[1687]=rom_data[12];
    rom_data[1688]=8'b10000110;
    rom_data[1689]=rom_data[12];
    rom_data[1690]=8'b10000110;
    rom_data[1691]=rom_data[12];
    rom_data[1692]=8'b10000110;
    rom_data[1693]=rom_data[12];
    rom_data[1694]=8'b10000110;
    rom_data[1695]=rom_data[12];
    rom_data[1696]=8'b10000110;
    rom_data[1697]=rom_data[12];
    rom_data[1698]=8'b10000101;
    rom_data[1699]=rom_data[12];
    rom_data[1700]=8'b10000101;
    rom_data[1701]=rom_data[12];
    rom_data[1702]=8'b10000101;
    rom_data[1703]=rom_data[12];
    rom_data[1704]=8'b10000101;
    rom_data[1705]=rom_data[12];
    rom_data[1706]=8'b10000101;
    rom_data[1707]=rom_data[12];
    rom_data[1708]=8'b10000101;
    rom_data[1709]=rom_data[12];
    rom_data[1710]=8'b10000101;
    rom_data[1711]=rom_data[12];
    rom_data[1712]=8'b10000101;
    rom_data[1713]=rom_data[12];
    rom_data[1714]=8'b10000100;
    rom_data[1715]=rom_data[12];
    rom_data[1716]=8'b10000100;
    rom_data[1717]=rom_data[12];
    rom_data[1718]=8'b10000100;
    rom_data[1719]=rom_data[12];
    rom_data[1720]=8'b10000100;
    rom_data[1721]=rom_data[12];
    rom_data[1722]=8'b10000100;
    rom_data[1723]=rom_data[12];
    rom_data[1724]=8'b10000100;
    rom_data[1725]=rom_data[12];
    rom_data[1726]=8'b10000100;
    rom_data[1727]=rom_data[12];
    rom_data[1728]=8'b10000011;
    rom_data[1729]=rom_data[12];
    rom_data[1730]=8'b10000011;
    rom_data[1731]=rom_data[12];
    rom_data[1732]=8'b10000011;
    rom_data[1733]=rom_data[12];
    rom_data[1734]=8'b10000011;
    rom_data[1735]=rom_data[12];
    rom_data[1736]=8'b10000011;
    rom_data[1737]=rom_data[12];
    rom_data[1738]=8'b10000011;
    rom_data[1739]=rom_data[12];
    rom_data[1740]=8'b10000011;
    rom_data[1741]=rom_data[12];
    rom_data[1742]=8'b10000011;
    rom_data[1743]=rom_data[12];
    rom_data[1744]=8'b10000010;
    rom_data[1745]=rom_data[12];
    rom_data[1746]=8'b10000010;
    rom_data[1747]=rom_data[12];
    rom_data[1748]=8'b10000010;
    rom_data[1749]=rom_data[12];
    rom_data[1750]=8'b10000010;
    rom_data[1751]=rom_data[12];
    rom_data[1752]=8'b10000010;
    rom_data[1753]=rom_data[12];
    rom_data[1754]=8'b10000010;
    rom_data[1755]=rom_data[12];
    rom_data[1756]=8'b10000010;
    rom_data[1757]=rom_data[12];
    rom_data[1758]=8'b10000010;
    rom_data[1759]=rom_data[12];
    rom_data[1760]=8'b10000010;
    rom_data[1761]=rom_data[12];
    rom_data[1762]=8'b10000001;
    rom_data[1763]=rom_data[12];
    rom_data[1764]=8'b10000001;
    rom_data[1765]=rom_data[12];
    rom_data[1766]=8'b10000001;
    rom_data[1767]=rom_data[12];
    rom_data[1768]=8'b10000001;
    rom_data[1769]=rom_data[12];
    rom_data[1770]=8'b10000001;
    rom_data[1771]=rom_data[12];
    rom_data[1772]=8'b10000001;
    rom_data[1773]=rom_data[12];
    rom_data[1774]=8'b10000001;
    rom_data[1775]=rom_data[12];
    rom_data[1776]=8'b10000001;
    rom_data[1777]=rom_data[12];
    rom_data[1778]=8'b10000001;
    rom_data[1779]=rom_data[12];
    rom_data[1780]=8'b10000000;
    rom_data[1781]=rom_data[12];
    rom_data[1782]=8'b10000000;
    rom_data[1783]=rom_data[12];
    rom_data[1784]=8'b10000000;
    rom_data[1785]=rom_data[12];
    rom_data[1786]=8'b10000000;
    rom_data[1787]=rom_data[12];
    rom_data[1788]=8'b10000000;
    rom_data[1789]=rom_data[12];
    rom_data[1790]=8'b10000000;
    rom_data[1791]=rom_data[12];
    rom_data[1792]=8'b10000000;
    rom_data[1793]=rom_data[12];
    rom_data[1794]=8'b10000000;
    rom_data[1795]=rom_data[12];
    rom_data[1796]=8'b10000000;
    rom_data[1797]=rom_data[12];
    rom_data[1798]=8'b10000000;
    rom_data[1799]=rom_data[12];
    rom_data[1800]=8'b01111111;
    rom_data[1801]=rom_data[12];
    rom_data[1802]=8'b01111111;
    rom_data[1803]=rom_data[12];
    rom_data[1804]=8'b01111111;
    rom_data[1805]=rom_data[12];
    rom_data[1806]=8'b01111111;
    rom_data[1807]=rom_data[12];
    rom_data[1808]=8'b01111111;
    rom_data[1809]=rom_data[12];
    rom_data[1810]=8'b01111111;
    rom_data[1811]=rom_data[12];
    rom_data[1812]=8'b01111111;
    rom_data[1813]=rom_data[12];
    rom_data[1814]=8'b01111111;
    rom_data[1815]=rom_data[12];
    rom_data[1816]=8'b01111111;
    rom_data[1817]=rom_data[12];
    rom_data[1818]=8'b01111111;
    rom_data[1819]=rom_data[12];
    rom_data[1820]=8'b01111110;
    rom_data[1821]=rom_data[12];
    rom_data[1822]=8'b01111110;
    rom_data[1823]=rom_data[12];
    rom_data[1824]=8'b01111110;
    rom_data[1825]=rom_data[12];
    rom_data[1826]=8'b01111110;
    rom_data[1827]=rom_data[12];
    rom_data[1828]=8'b01111110;
    rom_data[1829]=rom_data[12];
    rom_data[1830]=8'b01111110;
    rom_data[1831]=rom_data[12];
    rom_data[1832]=8'b01111110;
    rom_data[1833]=rom_data[12];
    rom_data[1834]=8'b01111110;
    rom_data[1835]=rom_data[12];
    rom_data[1836]=8'b01111110;
    rom_data[1837]=rom_data[12];
    rom_data[1838]=8'b01111110;
    rom_data[1839]=rom_data[12];
    rom_data[1840]=8'b01111101;
    rom_data[1841]=rom_data[12];
    rom_data[1842]=8'b01111101;
    rom_data[1843]=rom_data[12];
    rom_data[1844]=8'b01111101;
    rom_data[1845]=rom_data[12];
    rom_data[1846]=8'b01111101;
    rom_data[1847]=rom_data[12];
    rom_data[1848]=8'b01111101;
    rom_data[1849]=rom_data[12];
    rom_data[1850]=8'b01111101;
    rom_data[1851]=rom_data[12];
    rom_data[1852]=8'b01111101;
    rom_data[1853]=rom_data[12];
    rom_data[1854]=8'b01111101;
    rom_data[1855]=rom_data[12];
    rom_data[1856]=8'b01111100;
    rom_data[1857]=rom_data[12];
    rom_data[1858]=8'b01111100;
    rom_data[1859]=rom_data[12];
    rom_data[1860]=8'b01111100;
    rom_data[1861]=rom_data[12];
    rom_data[1862]=8'b01111100;
    rom_data[1863]=rom_data[12];
    rom_data[1864]=8'b01111100;
    rom_data[1865]=rom_data[12];
    rom_data[1866]=8'b01111100;
    rom_data[1867]=rom_data[12];
    rom_data[1868]=8'b01111100;
    rom_data[1869]=rom_data[12];
    rom_data[1870]=8'b01111100;
    rom_data[1871]=rom_data[12];
    rom_data[1872]=8'b01111011;
    rom_data[1873]=rom_data[12];
    rom_data[1874]=8'b01111011;
    rom_data[1875]=rom_data[12];
    rom_data[1876]=8'b01111011;
    rom_data[1877]=rom_data[12];
    rom_data[1878]=8'b01111011;
    rom_data[1879]=rom_data[12];
    rom_data[1880]=8'b01111011;
    rom_data[1881]=rom_data[12];
    rom_data[1882]=8'b01111011;
    rom_data[1883]=rom_data[12];
    rom_data[1884]=8'b01111011;
    rom_data[1885]=rom_data[12];
    rom_data[1886]=8'b01111011;
    rom_data[1887]=rom_data[12];
    rom_data[1888]=8'b01111010;
    rom_data[1889]=rom_data[12];
    rom_data[1890]=8'b01111010;
    rom_data[1891]=rom_data[12];
    rom_data[1892]=8'b01111010;
    rom_data[1893]=rom_data[12];
    rom_data[1894]=8'b01111010;
    rom_data[1895]=rom_data[12];
    rom_data[1896]=8'b01111010;
    rom_data[1897]=rom_data[12];
    rom_data[1898]=8'b01111010;
    rom_data[1899]=rom_data[12];
    rom_data[1900]=8'b01111010;
    rom_data[1901]=rom_data[12];
    rom_data[1902]=8'b01111001;
    rom_data[1903]=rom_data[12];
    rom_data[1904]=8'b01111001;
    rom_data[1905]=rom_data[12];
    rom_data[1906]=8'b01111001;
    rom_data[1907]=rom_data[12];
    rom_data[1908]=8'b01111001;
    rom_data[1909]=rom_data[12];
    rom_data[1910]=8'b01111001;
    rom_data[1911]=rom_data[12];
    rom_data[1912]=8'b01111001;
    rom_data[1913]=rom_data[12];
    rom_data[1914]=8'b01111001;
    rom_data[1915]=rom_data[12];
    rom_data[1916]=8'b01111000;
    rom_data[1917]=rom_data[12];
    rom_data[1918]=8'b01111000;
    rom_data[1919]=rom_data[12];
    rom_data[1920]=8'b01111000;
    rom_data[1921]=rom_data[12];
    rom_data[1922]=8'b01111000;
    rom_data[1923]=rom_data[12];
    rom_data[1924]=8'b01111000;
    rom_data[1925]=rom_data[12];
    rom_data[1926]=8'b01111000;
    rom_data[1927]=rom_data[12];
    rom_data[1928]=8'b01111000;
    rom_data[1929]=rom_data[12];
    rom_data[1930]=8'b01111000;
    rom_data[1931]=rom_data[12];
    rom_data[1932]=8'b01111000;
    rom_data[1933]=rom_data[12];
    rom_data[1934]=8'b01110111;
    rom_data[1935]=rom_data[12];
    rom_data[1936]=8'b01110111;
    rom_data[1937]=rom_data[12];
    rom_data[1938]=8'b01110111;
    rom_data[1939]=rom_data[12];
    rom_data[1940]=8'b01110111;
    rom_data[1941]=rom_data[12];
    rom_data[1942]=8'b01110111;
    rom_data[1943]=rom_data[12];
    rom_data[1944]=8'b01110111;
    rom_data[1945]=rom_data[12];
    rom_data[1946]=8'b01110111;
    rom_data[1947]=rom_data[12];
    rom_data[1948]=8'b01110111;
    rom_data[1949]=rom_data[12];
    rom_data[1950]=8'b01110111;
    rom_data[1951]=rom_data[12];
    rom_data[1952]=8'b01110110;
    rom_data[1953]=rom_data[12];
    rom_data[1954]=8'b01110110;
    rom_data[1955]=rom_data[12];
    rom_data[1956]=8'b01110110;
    rom_data[1957]=rom_data[12];
    rom_data[1958]=8'b01110110;
    rom_data[1959]=rom_data[12];
    rom_data[1960]=8'b01110110;
    rom_data[1961]=rom_data[12];
    rom_data[1962]=8'b01110110;
    rom_data[1963]=rom_data[12];
    rom_data[1964]=8'b01110110;
    rom_data[1965]=rom_data[12];
    rom_data[1966]=8'b01110110;
    rom_data[1967]=rom_data[12];
    rom_data[1968]=8'b01110110;
    rom_data[1969]=rom_data[12];
    rom_data[1970]=8'b01110110;
    rom_data[1971]=rom_data[12];
    rom_data[1972]=8'b01110101;
    rom_data[1973]=rom_data[12];
    rom_data[1974]=8'b01110101;
    rom_data[1975]=rom_data[12];
    rom_data[1976]=8'b01110101;
    rom_data[1977]=rom_data[12];
    rom_data[1978]=8'b01110101;
    rom_data[1979]=rom_data[12];
    rom_data[1980]=8'b01110101;
    rom_data[1981]=rom_data[12];
    rom_data[1982]=8'b01110101;
    rom_data[1983]=rom_data[12];
    rom_data[1984]=8'b01110101;
    rom_data[1985]=rom_data[12];
    rom_data[1986]=8'b01110101;
    rom_data[1987]=rom_data[12];
    rom_data[1988]=8'b01110101;
    rom_data[1989]=rom_data[12];
    rom_data[1990]=8'b01110101;
    rom_data[1991]=rom_data[12];
    rom_data[1992]=8'b01110100;
    rom_data[1993]=rom_data[12];
    rom_data[1994]=8'b01110100;
    rom_data[1995]=rom_data[12];
    rom_data[1996]=8'b01110100;
    rom_data[1997]=rom_data[12];
    rom_data[1998]=8'b01110100;
    rom_data[1999]=rom_data[12];
    rom_data[2000]=8'b01110100;
    rom_data[2001]=rom_data[12];
    rom_data[2002]=8'b01110100;
    rom_data[2003]=rom_data[12];
    rom_data[2004]=8'b01110100;
    rom_data[2005]=rom_data[12];
    rom_data[2006]=8'b01110100;
    rom_data[2007]=rom_data[12];
    rom_data[2008]=8'b01110100;
    rom_data[2009]=rom_data[12];
    rom_data[2010]=8'b01110100;
    rom_data[2011]=rom_data[12];
    rom_data[2012]=8'b01110011;
    rom_data[2013]=rom_data[12];
    rom_data[2014]=8'b01110011;
    rom_data[2015]=rom_data[12];
    rom_data[2016]=8'b01110011;
    rom_data[2017]=rom_data[12];
    rom_data[2018]=8'b01110011;
    rom_data[2019]=rom_data[12];
    rom_data[2020]=8'b01110011;
    rom_data[2021]=rom_data[12];
    rom_data[2022]=8'b01110011;
    rom_data[2023]=rom_data[12];
    rom_data[2024]=8'b01110011;
    rom_data[2025]=rom_data[12];
    rom_data[2026]=8'b01110011;
    rom_data[2027]=rom_data[12];
    rom_data[2028]=8'b01110011;
    rom_data[2029]=rom_data[12];
    rom_data[2030]=8'b01110010;
    rom_data[2031]=rom_data[12];
    rom_data[2032]=8'b01110010;
    rom_data[2033]=rom_data[12];
    rom_data[2034]=8'b01110010;
    rom_data[2035]=rom_data[12];
    rom_data[2036]=8'b01110010;
    rom_data[2037]=rom_data[12];
    rom_data[2038]=8'b01110010;
    rom_data[2039]=rom_data[12];
    rom_data[2040]=8'b01110010;
    rom_data[2041]=rom_data[12];
    rom_data[2042]=8'b01110010;
    rom_data[2043]=rom_data[12];
    rom_data[2044]=8'b01110010;
    rom_data[2045]=rom_data[12];
    rom_data[2046]=8'b01110001;
    rom_data[2047]=rom_data[12];
    rom_data[2048]=8'b01110001;
    rom_data[2049]=rom_data[12];
    rom_data[2050]=8'b01110001;
    rom_data[2051]=rom_data[12];
    rom_data[2052]=8'b01110001;
    rom_data[2053]=rom_data[12];
    rom_data[2054]=8'b01110001;
    rom_data[2055]=rom_data[12];
    rom_data[2056]=8'b01110001;
    rom_data[2057]=rom_data[12];
    rom_data[2058]=8'b01110001;
    rom_data[2059]=rom_data[12];
    rom_data[2060]=8'b01110000;
    rom_data[2061]=rom_data[12];
    rom_data[2062]=8'b01110000;
    rom_data[2063]=rom_data[12];
    rom_data[2064]=8'b01110000;
    rom_data[2065]=rom_data[12];
    rom_data[2066]=8'b01110000;
    rom_data[2067]=rom_data[12];
    rom_data[2068]=8'b01110000;
    rom_data[2069]=rom_data[12];
    rom_data[2070]=8'b01110000;
    rom_data[2071]=rom_data[12];
    rom_data[2072]=8'b01110000;
    rom_data[2073]=rom_data[12];
    rom_data[2074]=8'b01110000;
    rom_data[2075]=rom_data[12];
    rom_data[2076]=8'b01101111;
    rom_data[2077]=rom_data[12];
    rom_data[2078]=8'b01101111;
    rom_data[2079]=rom_data[12];
    rom_data[2080]=8'b01101111;
    rom_data[2081]=rom_data[12];
    rom_data[2082]=8'b01101111;
    rom_data[2083]=rom_data[12];
    rom_data[2084]=8'b01101111;
    rom_data[2085]=rom_data[12];
    rom_data[2086]=8'b01101111;
    rom_data[2087]=rom_data[12];
    rom_data[2088]=8'b01101111;
    rom_data[2089]=rom_data[12];
    rom_data[2090]=8'b01101110;
    rom_data[2091]=rom_data[12];
    rom_data[2092]=8'b01101110;
    rom_data[2093]=rom_data[12];
    rom_data[2094]=8'b01101110;
    rom_data[2095]=rom_data[12];
    rom_data[2096]=8'b01101110;
    rom_data[2097]=rom_data[12];
    rom_data[2098]=8'b01101110;
    rom_data[2099]=rom_data[12];
    rom_data[2100]=8'b01101110;
    rom_data[2101]=rom_data[12];
    rom_data[2102]=8'b01101110;
    rom_data[2103]=rom_data[12];
    rom_data[2104]=8'b01101110;
    rom_data[2105]=rom_data[12];
    rom_data[2106]=8'b01101101;
    rom_data[2107]=rom_data[12];
    rom_data[2108]=8'b01101101;
    rom_data[2109]=rom_data[12];
    rom_data[2110]=8'b01101101;
    rom_data[2111]=rom_data[12];
    rom_data[2112]=8'b01101101;
    rom_data[2113]=rom_data[12];
    rom_data[2114]=8'b01101101;
    rom_data[2115]=rom_data[12];
    rom_data[2116]=8'b01101101;
    rom_data[2117]=rom_data[12];
    rom_data[2118]=8'b01101101;
    rom_data[2119]=rom_data[12];
    rom_data[2120]=8'b01101101;
    rom_data[2121]=rom_data[12];
    rom_data[2122]=8'b01101101;
    rom_data[2123]=rom_data[12];
    rom_data[2124]=8'b01101100;
    rom_data[2125]=rom_data[12];
    rom_data[2126]=8'b01101100;
    rom_data[2127]=rom_data[12];
    rom_data[2128]=8'b01101100;
    rom_data[2129]=rom_data[12];
    rom_data[2130]=8'b01101100;
    rom_data[2131]=rom_data[12];
    rom_data[2132]=8'b01101100;
    rom_data[2133]=rom_data[12];
    rom_data[2134]=8'b01101100;
    rom_data[2135]=rom_data[12];
    rom_data[2136]=8'b01101100;
    rom_data[2137]=rom_data[12];
    rom_data[2138]=8'b01101100;
    rom_data[2139]=rom_data[12];
    rom_data[2140]=8'b01101100;
    rom_data[2141]=rom_data[12];
    rom_data[2142]=8'b01101100;
    rom_data[2143]=rom_data[12];
    rom_data[2144]=8'b01101011;
    rom_data[2145]=rom_data[12];
    rom_data[2146]=8'b01101011;
    rom_data[2147]=rom_data[12];
    rom_data[2148]=8'b01101011;
    rom_data[2149]=rom_data[12];
    rom_data[2150]=8'b01101011;
    rom_data[2151]=rom_data[12];
    rom_data[2152]=8'b01101011;
    rom_data[2153]=rom_data[12];
    rom_data[2154]=8'b01101011;
    rom_data[2155]=rom_data[12];
    rom_data[2156]=8'b01101011;
    rom_data[2157]=rom_data[12];
    rom_data[2158]=8'b01101011;
    rom_data[2159]=rom_data[12];
    rom_data[2160]=8'b01101011;
    rom_data[2161]=rom_data[12];
    rom_data[2162]=8'b01101011;
    rom_data[2163]=rom_data[12];
    rom_data[2164]=8'b01101010;
    rom_data[2165]=rom_data[12];
    rom_data[2166]=8'b01101010;
    rom_data[2167]=rom_data[12];
    rom_data[2168]=8'b01101010;
    rom_data[2169]=rom_data[12];
    rom_data[2170]=8'b01101010;
    rom_data[2171]=rom_data[12];
    rom_data[2172]=8'b01101010;
    rom_data[2173]=rom_data[12];
    rom_data[2174]=8'b01101010;
    rom_data[2175]=rom_data[12];
    rom_data[2176]=8'b01101010;
    rom_data[2177]=rom_data[12];
    rom_data[2178]=8'b01101010;
    rom_data[2179]=rom_data[12];
    rom_data[2180]=8'b01101010;
    rom_data[2181]=rom_data[12];
    rom_data[2182]=8'b01101001;
    rom_data[2183]=rom_data[12];
    rom_data[2184]=8'b01101001;
    rom_data[2185]=rom_data[12];
    rom_data[2186]=8'b01101001;
    rom_data[2187]=rom_data[12];
    rom_data[2188]=8'b01101001;
    rom_data[2189]=rom_data[12];
    rom_data[2190]=8'b01101001;
    rom_data[2191]=rom_data[12];
    rom_data[2192]=8'b01101001;
    rom_data[2193]=rom_data[12];
    rom_data[2194]=8'b01101001;
    rom_data[2195]=rom_data[12];
    rom_data[2196]=8'b01101001;
    rom_data[2197]=rom_data[12];
    rom_data[2198]=8'b01101001;
    rom_data[2199]=rom_data[12];
    rom_data[2200]=8'b01101001;
    rom_data[2201]=rom_data[12];
    rom_data[2202]=8'b01101000;
    rom_data[2203]=rom_data[12];
    rom_data[2204]=8'b01101000;
    rom_data[2205]=rom_data[12];
    rom_data[2206]=8'b01101000;
    rom_data[2207]=rom_data[12];
    rom_data[2208]=8'b01101000;
    rom_data[2209]=rom_data[12];
    rom_data[2210]=8'b01101000;
    rom_data[2211]=rom_data[12];
    rom_data[2212]=8'b01101000;
    rom_data[2213]=rom_data[12];
    rom_data[2214]=8'b01101000;
    rom_data[2215]=rom_data[12];
    rom_data[2216]=8'b01101000;
    rom_data[2217]=rom_data[12];
    rom_data[2218]=8'b01101000;
    rom_data[2219]=rom_data[12];
    rom_data[2220]=8'b01100111;
    rom_data[2221]=rom_data[12];
    rom_data[2222]=8'b01100111;
    rom_data[2223]=rom_data[12];
    rom_data[2224]=8'b01100111;
    rom_data[2225]=rom_data[12];
    rom_data[2226]=8'b01100111;
    rom_data[2227]=rom_data[12];
    rom_data[2228]=8'b01100111;
    rom_data[2229]=rom_data[12];
    rom_data[2230]=8'b01100111;
    rom_data[2231]=rom_data[12];
    rom_data[2232]=8'b01100111;
    rom_data[2233]=rom_data[12];
    rom_data[2234]=8'b01100110;
    rom_data[2235]=rom_data[12];
    rom_data[2236]=8'b01100110;
    rom_data[2237]=rom_data[12];
    rom_data[2238]=8'b01100110;
    rom_data[2239]=rom_data[12];
    rom_data[2240]=8'b01100110;
    rom_data[2241]=rom_data[12];
    rom_data[2242]=8'b01100110;
    rom_data[2243]=rom_data[12];
    rom_data[2244]=8'b01100110;
    rom_data[2245]=rom_data[12];
    rom_data[2246]=8'b01100110;
    rom_data[2247]=rom_data[12];
    rom_data[2248]=8'b01100110;
    rom_data[2249]=rom_data[12];
    rom_data[2250]=8'b01100101;
    rom_data[2251]=rom_data[12];
    rom_data[2252]=8'b01100101;
    rom_data[2253]=rom_data[12];
    rom_data[2254]=8'b01100101;
    rom_data[2255]=rom_data[12];
    rom_data[2256]=8'b01100101;
    rom_data[2257]=rom_data[12];
    rom_data[2258]=8'b01100101;
    rom_data[2259]=rom_data[12];
    rom_data[2260]=8'b01100101;
    rom_data[2261]=rom_data[12];
    rom_data[2262]=8'b01100101;
    rom_data[2263]=rom_data[12];
    rom_data[2264]=8'b01100100;
    rom_data[2265]=rom_data[12];
    rom_data[2266]=8'b01100100;
    rom_data[2267]=rom_data[12];
    rom_data[2268]=8'b01100100;
    rom_data[2269]=rom_data[12];
    rom_data[2270]=8'b01100100;
    rom_data[2271]=rom_data[12];
    rom_data[2272]=8'b01100100;
    rom_data[2273]=rom_data[12];
    rom_data[2274]=8'b01100100;
    rom_data[2275]=rom_data[12];
    rom_data[2276]=8'b01100100;
    rom_data[2277]=rom_data[12];
    rom_data[2278]=8'b01100011;
    rom_data[2279]=rom_data[12];
    rom_data[2280]=8'b01100011;
    rom_data[2281]=rom_data[12];
    rom_data[2282]=8'b01100011;
    rom_data[2283]=rom_data[12];
    rom_data[2284]=8'b01100011;
    rom_data[2285]=rom_data[12];
    rom_data[2286]=8'b01100011;
    rom_data[2287]=rom_data[12];
    rom_data[2288]=8'b01100011;
    rom_data[2289]=rom_data[12];
    rom_data[2290]=8'b01100011;
    rom_data[2291]=rom_data[12];
    rom_data[2292]=8'b01100011;
    rom_data[2293]=rom_data[12];
    rom_data[2294]=8'b01100011;
    rom_data[2295]=rom_data[12];
    rom_data[2296]=8'b01100010;
    rom_data[2297]=rom_data[12];
    rom_data[2298]=8'b01100010;
    rom_data[2299]=rom_data[12];
    rom_data[2300]=8'b01100010;
    rom_data[2301]=rom_data[12];
    rom_data[2302]=8'b01100010;
    rom_data[2303]=rom_data[12];
    rom_data[2304]=8'b01100010;
    rom_data[2305]=rom_data[12];
    rom_data[2306]=8'b01100010;
    rom_data[2307]=rom_data[12];
    rom_data[2308]=8'b01100010;
    rom_data[2309]=rom_data[12];
    rom_data[2310]=8'b01100010;
    rom_data[2311]=rom_data[12];
    rom_data[2312]=8'b01100010;
    rom_data[2313]=rom_data[12];
    rom_data[2314]=8'b01100001;
    rom_data[2315]=rom_data[12];
    rom_data[2316]=8'b01100001;
    rom_data[2317]=rom_data[12];
    rom_data[2318]=8'b01100001;
    rom_data[2319]=rom_data[12];
    rom_data[2320]=8'b01100001;
    rom_data[2321]=rom_data[12];
    rom_data[2322]=8'b01100001;
    rom_data[2323]=rom_data[12];
    rom_data[2324]=8'b01100001;
    rom_data[2325]=rom_data[12];
    rom_data[2326]=8'b01100001;
    rom_data[2327]=rom_data[12];
    rom_data[2328]=8'b01100001;
    rom_data[2329]=rom_data[12];
    rom_data[2330]=8'b01100001;
    rom_data[2331]=rom_data[12];
    rom_data[2332]=8'b01100001;
    rom_data[2333]=rom_data[12];
    rom_data[2334]=8'b01100000;
    rom_data[2335]=rom_data[12];
    rom_data[2336]=8'b01100000;
    rom_data[2337]=rom_data[12];
    rom_data[2338]=8'b01100000;
    rom_data[2339]=rom_data[12];
    rom_data[2340]=8'b01100000;
    rom_data[2341]=rom_data[12];
    rom_data[2342]=8'b01100000;
    rom_data[2343]=rom_data[12];
    rom_data[2344]=8'b01100000;
    rom_data[2345]=rom_data[12];
    rom_data[2346]=8'b01100000;
    rom_data[2347]=rom_data[12];
    rom_data[2348]=8'b01100000;
    rom_data[2349]=rom_data[12];
    rom_data[2350]=8'b01100000;
    rom_data[2351]=rom_data[12];
    rom_data[2352]=8'b01100000;
    rom_data[2353]=rom_data[12];
    rom_data[2354]=8'b01011111;
    rom_data[2355]=rom_data[12];
    rom_data[2356]=8'b01011111;
    rom_data[2357]=rom_data[12];
    rom_data[2358]=8'b01011111;
    rom_data[2359]=rom_data[12];
    rom_data[2360]=8'b01011111;
    rom_data[2361]=rom_data[12];
    rom_data[2362]=8'b01011111;
    rom_data[2363]=rom_data[12];
    rom_data[2364]=8'b01011111;
    rom_data[2365]=rom_data[12];
    rom_data[2366]=8'b01011111;
    rom_data[2367]=rom_data[12];
    rom_data[2368]=8'b01011111;
    rom_data[2369]=rom_data[12];
    rom_data[2370]=8'b01011111;
    rom_data[2371]=rom_data[12];
    rom_data[2372]=8'b01011111;
    rom_data[2373]=rom_data[12];
    rom_data[2374]=8'b01011110;
    rom_data[2375]=rom_data[12];
    rom_data[2376]=8'b01011110;
    rom_data[2377]=rom_data[12];
    rom_data[2378]=8'b01011110;
    rom_data[2379]=rom_data[12];
    rom_data[2380]=8'b01011110;
    rom_data[2381]=rom_data[12];
    rom_data[2382]=8'b01011110;
    rom_data[2383]=rom_data[12];
    rom_data[2384]=8'b01011110;
    rom_data[2385]=rom_data[12];
    rom_data[2386]=8'b01011110;
    rom_data[2387]=rom_data[12];
    rom_data[2388]=8'b01011110;
    rom_data[2389]=rom_data[12];
    rom_data[2390]=8'b01011110;
    rom_data[2391]=rom_data[12];
    rom_data[2392]=8'b01011101;
    rom_data[2393]=rom_data[12];
    rom_data[2394]=8'b01011101;
    rom_data[2395]=rom_data[12];
    rom_data[2396]=8'b01011101;
    rom_data[2397]=rom_data[12];
    rom_data[2398]=8'b01011101;
    rom_data[2399]=rom_data[12];
    rom_data[2400]=8'b01011101;
    rom_data[2401]=rom_data[12];
    rom_data[2402]=8'b01011101;
    rom_data[2403]=rom_data[12];
    rom_data[2404]=8'b01011101;
    rom_data[2405]=rom_data[12];
    rom_data[2406]=8'b01011101;
    rom_data[2407]=rom_data[12];
    rom_data[2408]=8'b01011100;
    rom_data[2409]=rom_data[12];
    rom_data[2410]=8'b01011100;
    rom_data[2411]=rom_data[12];
    rom_data[2412]=8'b01011100;
    rom_data[2413]=rom_data[12];
    rom_data[2414]=8'b01011100;
    rom_data[2415]=rom_data[12];
    rom_data[2416]=8'b01011100;
    rom_data[2417]=rom_data[12];
    rom_data[2418]=8'b01011100;
    rom_data[2419]=rom_data[12];
    rom_data[2420]=8'b01011100;
    rom_data[2421]=rom_data[12];
    rom_data[2422]=8'b01011011;
    rom_data[2423]=rom_data[12];
    rom_data[2424]=8'b01011011;
    rom_data[2425]=rom_data[12];
    rom_data[2426]=8'b01011011;
    rom_data[2427]=rom_data[12];
    rom_data[2428]=8'b01011011;
    rom_data[2429]=rom_data[12];
    rom_data[2430]=8'b01011011;
    rom_data[2431]=rom_data[12];
    rom_data[2432]=8'b01011011;
    rom_data[2433]=rom_data[12];
    rom_data[2434]=8'b01011011;
    rom_data[2435]=rom_data[12];
    rom_data[2436]=8'b01011011;
    rom_data[2437]=rom_data[12];
    rom_data[2438]=8'b01011010;
    rom_data[2439]=rom_data[12];
    rom_data[2440]=8'b01011010;
    rom_data[2441]=rom_data[12];
    rom_data[2442]=8'b01011010;
    rom_data[2443]=rom_data[12];
    rom_data[2444]=8'b01011010;
    rom_data[2445]=rom_data[12];
    rom_data[2446]=8'b01011010;
    rom_data[2447]=rom_data[12];
    rom_data[2448]=8'b01011010;
    rom_data[2449]=rom_data[12];
    rom_data[2450]=8'b01011010;
    rom_data[2451]=rom_data[12];
    rom_data[2452]=8'b01011001;
    rom_data[2453]=rom_data[12];
    rom_data[2454]=8'b01011001;
    rom_data[2455]=rom_data[12];
    rom_data[2456]=8'b01011001;
    rom_data[2457]=rom_data[12];
    rom_data[2458]=8'b01011001;
    rom_data[2459]=rom_data[12];
    rom_data[2460]=8'b01011001;
    rom_data[2461]=rom_data[12];
    rom_data[2462]=8'b01011001;
    rom_data[2463]=rom_data[12];
    rom_data[2464]=8'b01011001;
    rom_data[2465]=rom_data[12];
    rom_data[2466]=8'b01011001;
    rom_data[2467]=rom_data[12];
    rom_data[2468]=8'b01011000;
    rom_data[2469]=rom_data[12];
    rom_data[2470]=8'b01011000;
    rom_data[2471]=rom_data[12];
    rom_data[2472]=8'b01011000;
    rom_data[2473]=rom_data[12];
    rom_data[2474]=8'b01011000;
    rom_data[2475]=rom_data[12];
    rom_data[2476]=8'b01011000;
    rom_data[2477]=rom_data[12];
    rom_data[2478]=8'b01011000;
    rom_data[2479]=rom_data[12];
    rom_data[2480]=8'b01011000;
    rom_data[2481]=rom_data[12];
    rom_data[2482]=8'b01011000;
    rom_data[2483]=rom_data[12];
    rom_data[2484]=8'b01011000;
    rom_data[2485]=rom_data[12];
    rom_data[2486]=8'b01010111;
    rom_data[2487]=rom_data[12];
    rom_data[2488]=8'b01010111;
    rom_data[2489]=rom_data[12];
    rom_data[2490]=8'b01010111;
    rom_data[2491]=rom_data[12];
    rom_data[2492]=8'b01010111;
    rom_data[2493]=rom_data[12];
    rom_data[2494]=8'b01010111;
    rom_data[2495]=rom_data[12];
    rom_data[2496]=8'b01010111;
    rom_data[2497]=rom_data[12];
    rom_data[2498]=8'b01010111;
    rom_data[2499]=rom_data[12];
    rom_data[2500]=8'b01010111;
    rom_data[2501]=rom_data[12];
    rom_data[2502]=8'b01010111;
    rom_data[2503]=rom_data[12];
    rom_data[2504]=8'b01010111;
    rom_data[2505]=rom_data[12];
    rom_data[2506]=8'b01010110;
    rom_data[2507]=rom_data[12];
    rom_data[2508]=8'b01010110;
    rom_data[2509]=rom_data[12];
    rom_data[2510]=8'b01010110;
    rom_data[2511]=rom_data[12];
    rom_data[2512]=8'b01010110;
    rom_data[2513]=rom_data[12];
    rom_data[2514]=8'b01010110;
    rom_data[2515]=rom_data[12];
    rom_data[2516]=8'b01010110;
    rom_data[2517]=rom_data[12];
    rom_data[2518]=8'b01010110;
    rom_data[2519]=rom_data[12];
    rom_data[2520]=8'b01010110;
    rom_data[2521]=rom_data[12];
    rom_data[2522]=8'b01010110;
    rom_data[2523]=rom_data[12];
    rom_data[2524]=8'b01010110;
    rom_data[2525]=rom_data[12];
    rom_data[2526]=8'b01010101;
    rom_data[2527]=rom_data[12];
    rom_data[2528]=8'b01010101;
    rom_data[2529]=rom_data[12];
    rom_data[2530]=8'b01010101;
    rom_data[2531]=rom_data[12];
    rom_data[2532]=8'b01010101;
    rom_data[2533]=rom_data[12];
    rom_data[2534]=8'b01010101;
    rom_data[2535]=rom_data[12];
    rom_data[2536]=8'b01010101;
    rom_data[2537]=rom_data[12];
    rom_data[2538]=8'b01010101;
    rom_data[2539]=rom_data[12];
    rom_data[2540]=8'b01010101;
    rom_data[2541]=rom_data[12];
    rom_data[2542]=8'b01010101;
    rom_data[2543]=rom_data[12];
    rom_data[2544]=8'b01010101;
    rom_data[2545]=rom_data[12];
    rom_data[2546]=8'b01010100;
    rom_data[2547]=rom_data[12];
    rom_data[2548]=8'b01010100;
    rom_data[2549]=rom_data[12];
    rom_data[2550]=8'b01010100;
    rom_data[2551]=rom_data[12];
    rom_data[2552]=8'b01010100;
    rom_data[2553]=rom_data[12];
    rom_data[2554]=8'b01010100;
    rom_data[2555]=rom_data[12];
    rom_data[2556]=8'b01010100;
    rom_data[2557]=rom_data[12];
    rom_data[2558]=8'b01010100;
    rom_data[2559]=rom_data[12];
    rom_data[2560]=8'b01010100;
    rom_data[2561]=rom_data[12];
    rom_data[2562]=8'b01010100;
    rom_data[2563]=rom_data[12];
    rom_data[2564]=8'b01010011;
    rom_data[2565]=rom_data[12];
    rom_data[2566]=8'b01010011;
    rom_data[2567]=rom_data[12];
    rom_data[2568]=8'b01010011;
    rom_data[2569]=rom_data[12];
    rom_data[2570]=8'b01010011;
    rom_data[2571]=rom_data[12];
    rom_data[2572]=8'b01010011;
    rom_data[2573]=rom_data[12];
    rom_data[2574]=8'b01010011;
    rom_data[2575]=rom_data[12];
    rom_data[2576]=8'b01010011;
    rom_data[2577]=rom_data[12];
    rom_data[2578]=8'b01010011;
    rom_data[2579]=rom_data[12];
    rom_data[2580]=8'b01010011;
    rom_data[2581]=rom_data[12];
    rom_data[2582]=8'b01010010;
    rom_data[2583]=rom_data[12];
    rom_data[2584]=8'b01010010;
    rom_data[2585]=rom_data[12];
    rom_data[2586]=8'b01010010;
    rom_data[2587]=rom_data[12];
    rom_data[2588]=8'b01010010;
    rom_data[2589]=rom_data[12];
    rom_data[2590]=8'b01010010;
    rom_data[2591]=rom_data[12];
    rom_data[2592]=8'b01010010;
    rom_data[2593]=rom_data[12];
    rom_data[2594]=8'b01010010;
    rom_data[2595]=rom_data[12];
    rom_data[2596]=8'b01010001;
    rom_data[2597]=rom_data[12];
    rom_data[2598]=8'b01010001;
    rom_data[2599]=rom_data[12];
    rom_data[2600]=8'b01010001;
    rom_data[2601]=rom_data[12];
    rom_data[2602]=8'b01010001;
    rom_data[2603]=rom_data[12];
    rom_data[2604]=8'b01010001;
    rom_data[2605]=rom_data[12];
    rom_data[2606]=8'b01010001;
    rom_data[2607]=rom_data[12];
    rom_data[2608]=8'b01010001;
    rom_data[2609]=rom_data[12];
    rom_data[2610]=8'b01010001;
    rom_data[2611]=rom_data[12];
    rom_data[2612]=8'b01010000;
    rom_data[2613]=rom_data[12];
    rom_data[2614]=8'b01010000;
    rom_data[2615]=rom_data[12];
    rom_data[2616]=8'b01010000;
    rom_data[2617]=rom_data[12];
    rom_data[2618]=8'b01010000;
    rom_data[2619]=rom_data[12];
    rom_data[2620]=8'b01010000;
    rom_data[2621]=rom_data[12];
    rom_data[2622]=8'b01010000;
    rom_data[2623]=rom_data[12];
    rom_data[2624]=8'b01010000;
    rom_data[2625]=rom_data[12];
    rom_data[2626]=8'b01001111;
    rom_data[2627]=rom_data[12];
    rom_data[2628]=8'b01001111;
    rom_data[2629]=rom_data[12];
    rom_data[2630]=8'b01001111;
    rom_data[2631]=rom_data[12];
    rom_data[2632]=8'b01001111;
    rom_data[2633]=rom_data[12];
    rom_data[2634]=8'b01001111;
    rom_data[2635]=rom_data[12];
    rom_data[2636]=8'b01001111;
    rom_data[2637]=rom_data[12];
    rom_data[2638]=8'b01001111;
    rom_data[2639]=rom_data[12];
    rom_data[2640]=8'b01001111;
    rom_data[2641]=rom_data[12];
    rom_data[2642]=8'b01001110;
    rom_data[2643]=rom_data[12];
    rom_data[2644]=8'b01001110;
    rom_data[2645]=rom_data[12];
    rom_data[2646]=8'b01001110;
    rom_data[2647]=rom_data[12];
    rom_data[2648]=8'b01001110;
    rom_data[2649]=rom_data[12];
    rom_data[2650]=8'b01001110;
    rom_data[2651]=rom_data[12];
    rom_data[2652]=8'b01001110;
    rom_data[2653]=rom_data[12];
    rom_data[2654]=8'b01001110;
    rom_data[2655]=rom_data[12];
    rom_data[2656]=8'b01001110;
    rom_data[2657]=rom_data[12];
    rom_data[2658]=8'b01001101;
    rom_data[2659]=rom_data[12];
    rom_data[2660]=8'b01001101;
    rom_data[2661]=rom_data[12];
    rom_data[2662]=8'b01001101;
    rom_data[2663]=rom_data[12];
    rom_data[2664]=8'b01001101;
    rom_data[2665]=rom_data[12];
    rom_data[2666]=8'b01001101;
    rom_data[2667]=rom_data[12];
    rom_data[2668]=8'b01001101;
    rom_data[2669]=rom_data[12];
    rom_data[2670]=8'b01001101;
    rom_data[2671]=rom_data[12];
    rom_data[2672]=8'b01001101;
    rom_data[2673]=rom_data[12];
    rom_data[2674]=8'b01001101;
    rom_data[2675]=rom_data[12];
    rom_data[2676]=8'b01001101;
    rom_data[2677]=rom_data[12];
    rom_data[2678]=8'b01001100;
    rom_data[2679]=rom_data[12];
    rom_data[2680]=8'b01001100;
    rom_data[2681]=rom_data[12];
    rom_data[2682]=8'b01001100;
    rom_data[2683]=rom_data[12];
    rom_data[2684]=8'b01001100;
    rom_data[2685]=rom_data[12];
    rom_data[2686]=8'b01001100;
    rom_data[2687]=rom_data[12];
    rom_data[2688]=8'b01001100;
    rom_data[2689]=rom_data[12];
    rom_data[2690]=8'b01001100;
    rom_data[2691]=rom_data[12];
    rom_data[2692]=8'b01001100;
    rom_data[2693]=rom_data[12];
    rom_data[2694]=8'b01001100;
    rom_data[2695]=rom_data[12];
    rom_data[2696]=8'b01001100;
    rom_data[2697]=rom_data[12];
    rom_data[2698]=8'b01001011;
    rom_data[2699]=rom_data[12];
    rom_data[2700]=8'b01001011;
    rom_data[2701]=rom_data[12];
    rom_data[2702]=8'b01001011;
    rom_data[2703]=rom_data[12];
    rom_data[2704]=8'b01001011;
    rom_data[2705]=rom_data[12];
    rom_data[2706]=8'b01001011;
    rom_data[2707]=rom_data[12];
    rom_data[2708]=8'b01001011;
    rom_data[2709]=rom_data[12];
    rom_data[2710]=8'b01001011;
    rom_data[2711]=rom_data[12];
    rom_data[2712]=8'b01001011;
    rom_data[2713]=rom_data[12];
    rom_data[2714]=8'b01001011;
    rom_data[2715]=rom_data[12];
    rom_data[2716]=8'b01001011;
    rom_data[2717]=rom_data[12];
    rom_data[2718]=8'b01001010;
    rom_data[2719]=rom_data[12];
    rom_data[2720]=8'b01001010;
    rom_data[2721]=rom_data[12];
    rom_data[2722]=8'b01001010;
    rom_data[2723]=rom_data[12];
    rom_data[2724]=8'b01001010;
    rom_data[2725]=rom_data[12];
    rom_data[2726]=8'b01001010;
    rom_data[2727]=rom_data[12];
    rom_data[2728]=8'b01001010;
    rom_data[2729]=rom_data[12];
    rom_data[2730]=8'b01001010;
    rom_data[2731]=rom_data[12];
    rom_data[2732]=8'b01001010;
    rom_data[2733]=rom_data[12];
    rom_data[2734]=8'b01001010;
    rom_data[2735]=rom_data[12];
    rom_data[2736]=8'b01001001;
    rom_data[2737]=rom_data[12];
    rom_data[2738]=8'b01001001;
    rom_data[2739]=rom_data[12];
    rom_data[2740]=8'b01001001;
    rom_data[2741]=rom_data[12];
    rom_data[2742]=8'b01001001;
    rom_data[2743]=rom_data[12];
    rom_data[2744]=8'b01001001;
    rom_data[2745]=rom_data[12];
    rom_data[2746]=8'b01001001;
    rom_data[2747]=rom_data[12];
    rom_data[2748]=8'b01001001;
    rom_data[2749]=rom_data[12];
    rom_data[2750]=8'b01001001;
    rom_data[2751]=rom_data[12];
    rom_data[2752]=8'b01001001;
    rom_data[2753]=rom_data[12];
    rom_data[2754]=8'b01001000;
    rom_data[2755]=rom_data[12];
    rom_data[2756]=8'b01001000;
    rom_data[2757]=rom_data[12];
    rom_data[2758]=8'b01001000;
    rom_data[2759]=rom_data[12];
    rom_data[2760]=8'b01001000;
    rom_data[2761]=rom_data[12];
    rom_data[2762]=8'b01001000;
    rom_data[2763]=rom_data[12];
    rom_data[2764]=8'b01001000;
    rom_data[2765]=rom_data[12];
    rom_data[2766]=8'b01001000;
    rom_data[2767]=rom_data[12];
    rom_data[2768]=8'b01001000;
    rom_data[2769]=rom_data[12];
    rom_data[2770]=8'b01000111;
    rom_data[2771]=rom_data[12];
    rom_data[2772]=8'b01000111;
    rom_data[2773]=rom_data[12];
    rom_data[2774]=8'b01000111;
    rom_data[2775]=rom_data[12];
    rom_data[2776]=8'b01000111;
    rom_data[2777]=rom_data[12];
    rom_data[2778]=8'b01000111;
    rom_data[2779]=rom_data[12];
    rom_data[2780]=8'b01000111;
    rom_data[2781]=rom_data[12];
    rom_data[2782]=8'b01000111;
    rom_data[2783]=rom_data[12];
    rom_data[2784]=8'b01000111;
    rom_data[2785]=rom_data[12];
    rom_data[2786]=8'b01000110;
    rom_data[2787]=rom_data[12];
    rom_data[2788]=8'b01000110;
    rom_data[2789]=rom_data[12];
    rom_data[2790]=8'b01000110;
    rom_data[2791]=rom_data[12];
    rom_data[2792]=8'b01000110;
    rom_data[2793]=rom_data[12];
    rom_data[2794]=8'b01000110;
    rom_data[2795]=rom_data[12];
    rom_data[2796]=8'b01000110;
    rom_data[2797]=rom_data[12];
    rom_data[2798]=8'b01000110;
    rom_data[2799]=rom_data[12];
    rom_data[2800]=8'b01000101;
    rom_data[2801]=rom_data[12];
    rom_data[2802]=8'b01000101;
    rom_data[2803]=rom_data[12];
    rom_data[2804]=8'b01000101;
    rom_data[2805]=rom_data[12];
    rom_data[2806]=8'b01000101;
    rom_data[2807]=rom_data[12];
    rom_data[2808]=8'b01000101;
    rom_data[2809]=rom_data[12];
    rom_data[2810]=8'b01000101;
    rom_data[2811]=rom_data[12];
    rom_data[2812]=8'b01000101;
    rom_data[2813]=rom_data[12];
    rom_data[2814]=8'b01000100;
    rom_data[2815]=rom_data[12];
    rom_data[2816]=8'b01000100;
    rom_data[2817]=rom_data[12];
    rom_data[2818]=8'b01000100;
    rom_data[2819]=rom_data[12];
    rom_data[2820]=8'b01000100;
    rom_data[2821]=rom_data[12];
    rom_data[2822]=8'b01000100;
    rom_data[2823]=rom_data[12];
    rom_data[2824]=8'b01000100;
    rom_data[2825]=rom_data[12];
    rom_data[2826]=8'b01000100;
    rom_data[2827]=rom_data[12];
    rom_data[2828]=8'b01000100;
    rom_data[2829]=rom_data[12];
    rom_data[2830]=8'b01000011;
    rom_data[2831]=rom_data[12];
    rom_data[2832]=8'b01000011;
    rom_data[2833]=rom_data[12];
    rom_data[2834]=8'b01000011;
    rom_data[2835]=rom_data[12];
    rom_data[2836]=8'b01000011;
    rom_data[2837]=rom_data[12];
    rom_data[2838]=8'b01000011;
    rom_data[2839]=rom_data[12];
    rom_data[2840]=8'b01000011;
    rom_data[2841]=rom_data[12];
    rom_data[2842]=8'b01000011;
    rom_data[2843]=rom_data[12];
    rom_data[2844]=8'b01000011;
    rom_data[2845]=rom_data[12];
    rom_data[2846]=8'b01000011;
    rom_data[2847]=rom_data[12];
    rom_data[2848]=8'b01000011;
    rom_data[2849]=rom_data[12];
    rom_data[2850]=8'b01000010;
    rom_data[2851]=rom_data[12];
    rom_data[2852]=8'b01000010;
    rom_data[2853]=rom_data[12];
    rom_data[2854]=8'b01000010;
    rom_data[2855]=rom_data[12];
    rom_data[2856]=8'b01000010;
    rom_data[2857]=rom_data[12];
    rom_data[2858]=8'b01000010;
    rom_data[2859]=rom_data[12];
    rom_data[2860]=8'b01000010;
    rom_data[2861]=rom_data[12];
    rom_data[2862]=8'b01000010;
    rom_data[2863]=rom_data[12];
    rom_data[2864]=8'b01000010;
    rom_data[2865]=rom_data[12];
    rom_data[2866]=8'b01000010;
    rom_data[2867]=rom_data[12];
    rom_data[2868]=8'b01000001;
    rom_data[2869]=rom_data[12];
    rom_data[2870]=8'b01000001;
    rom_data[2871]=rom_data[12];
    rom_data[2872]=8'b01000001;
    rom_data[2873]=rom_data[12];
    rom_data[2874]=8'b01000001;
    rom_data[2875]=rom_data[12];
    rom_data[2876]=8'b01000001;
    rom_data[2877]=rom_data[12];
    rom_data[2878]=8'b01000001;
    rom_data[2879]=rom_data[12];
    rom_data[2880]=8'b01000001;
    rom_data[2881]=rom_data[12];
    rom_data[2882]=8'b01000001;
    rom_data[2883]=rom_data[12];
    rom_data[2884]=8'b01000001;
    rom_data[2885]=rom_data[12];
    rom_data[2886]=8'b01000001;
    rom_data[2887]=rom_data[12];
    rom_data[2888]=8'b01000000;
    rom_data[2889]=rom_data[12];
    rom_data[2890]=8'b01000000;
    rom_data[2891]=rom_data[12];
    rom_data[2892]=8'b01000000;
    rom_data[2893]=rom_data[12];
    rom_data[2894]=8'b01000000;
    rom_data[2895]=rom_data[12];
    rom_data[2896]=8'b01000000;
    rom_data[2897]=rom_data[12];
    rom_data[2898]=8'b01000000;
    rom_data[2899]=rom_data[12];
    rom_data[2900]=8'b01000000;
    rom_data[2901]=rom_data[12];
    rom_data[2902]=8'b01000000;
    rom_data[2903]=rom_data[12];
    rom_data[2904]=8'b01000000;
    rom_data[2905]=rom_data[12];
    rom_data[2906]=8'b01000000;
    rom_data[2907]=rom_data[12];
    rom_data[2908]=8'b00111111;
    rom_data[2909]=rom_data[12];
    rom_data[2910]=8'b00111111;
    rom_data[2911]=rom_data[12];
    rom_data[2912]=8'b00111111;
    rom_data[2913]=rom_data[12];
    rom_data[2914]=8'b00111111;
    rom_data[2915]=rom_data[12];
    rom_data[2916]=8'b00111111;
    rom_data[2917]=rom_data[12];
    rom_data[2918]=8'b00111111;
    rom_data[2919]=rom_data[12];
    rom_data[2920]=8'b00111111;
    rom_data[2921]=rom_data[12];
    rom_data[2922]=8'b00111111;
    rom_data[2923]=rom_data[12];
    rom_data[2924]=8'b00111111;
    rom_data[2925]=rom_data[12];
    rom_data[2926]=8'b00111110;
    rom_data[2927]=rom_data[12];
    rom_data[2928]=8'b00111110;
    rom_data[2929]=rom_data[12];
    rom_data[2930]=8'b00111110;
    rom_data[2931]=rom_data[12];
    rom_data[2932]=8'b00111110;
    rom_data[2933]=rom_data[12];
    rom_data[2934]=8'b00111110;
    rom_data[2935]=rom_data[12];
    rom_data[2936]=8'b00111110;
    rom_data[2937]=rom_data[12];
    rom_data[2938]=8'b00111110;
    rom_data[2939]=rom_data[12];
    rom_data[2940]=8'b00111110;
    rom_data[2941]=rom_data[12];
    rom_data[2942]=8'b00111110;
    rom_data[2943]=rom_data[12];
    rom_data[2944]=8'b00111101;
    rom_data[2945]=rom_data[12];
    rom_data[2946]=8'b00111101;
    rom_data[2947]=rom_data[12];
    rom_data[2948]=8'b00111101;
    rom_data[2949]=rom_data[12];
    rom_data[2950]=8'b00111101;
    rom_data[2951]=rom_data[12];
    rom_data[2952]=8'b00111101;
    rom_data[2953]=rom_data[12];
    rom_data[2954]=8'b00111101;
    rom_data[2955]=rom_data[12];
    rom_data[2956]=8'b00111101;
    rom_data[2957]=rom_data[12];
    rom_data[2958]=8'b00111100;
    rom_data[2959]=rom_data[12];
    rom_data[2960]=8'b00111100;
    rom_data[2961]=rom_data[12];
    rom_data[2962]=8'b00111100;
    rom_data[2963]=rom_data[12];
    rom_data[2964]=8'b00111100;
    rom_data[2965]=rom_data[12];
    rom_data[2966]=8'b00111100;
    rom_data[2967]=rom_data[12];
    rom_data[2968]=8'b00111100;
    rom_data[2969]=rom_data[12];
    rom_data[2970]=8'b00111100;
    rom_data[2971]=rom_data[12];
    rom_data[2972]=8'b00111100;
    rom_data[2973]=rom_data[12];
    rom_data[2974]=8'b00111011;
    rom_data[2975]=rom_data[12];
    rom_data[2976]=8'b00111011;
    rom_data[2977]=rom_data[12];
    rom_data[2978]=8'b00111011;
    rom_data[2979]=rom_data[12];
    rom_data[2980]=8'b00111011;
    rom_data[2981]=rom_data[12];
    rom_data[2982]=8'b00111011;
    rom_data[2983]=rom_data[12];
    rom_data[2984]=8'b00111011;
    rom_data[2985]=rom_data[12];
    rom_data[2986]=8'b00111011;
    rom_data[2987]=rom_data[12];
    rom_data[2988]=8'b00111010;
    rom_data[2989]=rom_data[12];
    rom_data[2990]=8'b00111010;
    rom_data[2991]=rom_data[12];
    rom_data[2992]=8'b00111010;
    rom_data[2993]=rom_data[12];
    rom_data[2994]=8'b00111010;
    rom_data[2995]=rom_data[12];
    rom_data[2996]=8'b00111010;
    rom_data[2997]=rom_data[12];
    rom_data[2998]=8'b00111010;
    rom_data[2999]=rom_data[12];
    rom_data[3000]=8'b00111010;
    rom_data[3001]=rom_data[12];
    rom_data[3002]=8'b00111010;
    rom_data[3003]=rom_data[12];
    rom_data[3004]=8'b00111001;
    rom_data[3005]=rom_data[12];
    rom_data[3006]=8'b00111001;
    rom_data[3007]=rom_data[12];
    rom_data[3008]=8'b00111001;
    rom_data[3009]=rom_data[12];
    rom_data[3010]=8'b00111001;
    rom_data[3011]=rom_data[12];
    rom_data[3012]=8'b00111001;
    rom_data[3013]=rom_data[12];
    rom_data[3014]=8'b00111001;
    rom_data[3015]=rom_data[12];
    rom_data[3016]=8'b00111001;
    rom_data[3017]=rom_data[12];
    rom_data[3018]=8'b00111001;
    rom_data[3019]=rom_data[12];
    rom_data[3020]=8'b00111001;
    rom_data[3021]=rom_data[12];
    rom_data[3022]=8'b00111000;
    rom_data[3023]=rom_data[12];
    rom_data[3024]=8'b00111000;
    rom_data[3025]=rom_data[12];
    rom_data[3026]=8'b00111000;
    rom_data[3027]=rom_data[12];
    rom_data[3028]=8'b00111000;
    rom_data[3029]=rom_data[12];
    rom_data[3030]=8'b00111000;
    rom_data[3031]=rom_data[12];
    rom_data[3032]=8'b00111000;
    rom_data[3033]=rom_data[12];
    rom_data[3034]=8'b00111000;
    rom_data[3035]=rom_data[12];
    rom_data[3036]=8'b00111000;
    rom_data[3037]=rom_data[12];
    rom_data[3038]=8'b00111000;
    rom_data[3039]=rom_data[12];
    rom_data[3040]=8'b00110111;
    rom_data[3041]=rom_data[12];
    rom_data[3042]=8'b00110111;
    rom_data[3043]=rom_data[12];
    rom_data[3044]=8'b00110111;
    rom_data[3045]=rom_data[12];
    rom_data[3046]=8'b00110111;
    rom_data[3047]=rom_data[12];
    rom_data[3048]=8'b00110111;
    rom_data[3049]=rom_data[12];
    rom_data[3050]=8'b00110111;
    rom_data[3051]=rom_data[12];
    rom_data[3052]=8'b00110111;
    rom_data[3053]=rom_data[12];
    rom_data[3054]=8'b00110111;
    rom_data[3055]=rom_data[12];
    rom_data[3056]=8'b00110111;
    rom_data[3057]=rom_data[12];
    rom_data[3058]=8'b00110111;
    rom_data[3059]=rom_data[12];
    rom_data[3060]=8'b00110110;
    rom_data[3061]=rom_data[12];
    rom_data[3062]=8'b00110110;
    rom_data[3063]=rom_data[12];
    rom_data[3064]=8'b00110110;
    rom_data[3065]=rom_data[12];
    rom_data[3066]=8'b00110110;
    rom_data[3067]=rom_data[12];
    rom_data[3068]=8'b00110110;
    rom_data[3069]=rom_data[12];
    rom_data[3070]=8'b00110110;
    rom_data[3071]=rom_data[12];
    rom_data[3072]=8'b00110110;
    rom_data[3073]=rom_data[12];
    rom_data[3074]=8'b00110110;
    rom_data[3075]=rom_data[12];
    rom_data[3076]=8'b00110110;
    rom_data[3077]=rom_data[12];
    rom_data[3078]=8'b00110110;
    rom_data[3079]=rom_data[12];
    rom_data[3080]=8'b00110101;
    rom_data[3081]=rom_data[12];
    rom_data[3082]=8'b00110101;
    rom_data[3083]=rom_data[12];
    rom_data[3084]=8'b00110101;
    rom_data[3085]=rom_data[12];
    rom_data[3086]=8'b00110101;
    rom_data[3087]=rom_data[12];
    rom_data[3088]=8'b00110101;
    rom_data[3089]=rom_data[12];
    rom_data[3090]=8'b00110101;
    rom_data[3091]=rom_data[12];
    rom_data[3092]=8'b00110101;
    rom_data[3093]=rom_data[12];
    rom_data[3094]=8'b00110101;
    rom_data[3095]=rom_data[12];
    rom_data[3096]=8'b00110101;
    rom_data[3097]=rom_data[12];
    rom_data[3098]=8'b00110101;
    rom_data[3099]=rom_data[12];
    rom_data[3100]=8'b00110100;
    rom_data[3101]=rom_data[12];
    rom_data[3102]=8'b00110100;
    rom_data[3103]=rom_data[12];
    rom_data[3104]=8'b00110100;
    rom_data[3105]=rom_data[12];
    rom_data[3106]=8'b00110100;
    rom_data[3107]=rom_data[12];
    rom_data[3108]=8'b00110100;
    rom_data[3109]=rom_data[12];
    rom_data[3110]=8'b00110100;
    rom_data[3111]=rom_data[12];
    rom_data[3112]=8'b00110100;
    rom_data[3113]=rom_data[12];
    rom_data[3114]=8'b00110100;
    rom_data[3115]=rom_data[12];
    rom_data[3116]=8'b00110011;
    rom_data[3117]=rom_data[12];
    rom_data[3118]=8'b00110011;
    rom_data[3119]=rom_data[12];
    rom_data[3120]=8'b00110011;
    rom_data[3121]=rom_data[12];
    rom_data[3122]=8'b00110011;
    rom_data[3123]=rom_data[12];
    rom_data[3124]=8'b00110011;
    rom_data[3125]=rom_data[12];
    rom_data[3126]=8'b00110011;
    rom_data[3127]=rom_data[12];
    rom_data[3128]=8'b00110011;
    rom_data[3129]=rom_data[12];
    rom_data[3130]=8'b00110011;
    rom_data[3131]=rom_data[12];
    rom_data[3132]=8'b00110010;
    rom_data[3133]=rom_data[12];
    rom_data[3134]=8'b00110010;
    rom_data[3135]=rom_data[12];
    rom_data[3136]=8'b00110010;
    rom_data[3137]=rom_data[12];
    rom_data[3138]=8'b00110010;
    rom_data[3139]=rom_data[12];
    rom_data[3140]=8'b00110010;
    rom_data[3141]=rom_data[12];
    rom_data[3142]=8'b00110010;
    rom_data[3143]=rom_data[12];
    rom_data[3144]=8'b00110010;
    rom_data[3145]=rom_data[12];
    rom_data[3146]=8'b00110010;
    rom_data[3147]=rom_data[12];
    rom_data[3148]=8'b00110001;
    rom_data[3149]=rom_data[12];
    rom_data[3150]=8'b00110001;
    rom_data[3151]=rom_data[12];
    rom_data[3152]=8'b00110001;
    rom_data[3153]=rom_data[12];
    rom_data[3154]=8'b00110001;
    rom_data[3155]=rom_data[12];
    rom_data[3156]=8'b00110001;
    rom_data[3157]=rom_data[12];
    rom_data[3158]=8'b00110001;
    rom_data[3159]=rom_data[12];
    rom_data[3160]=8'b00110001;
    rom_data[3161]=rom_data[12];
    rom_data[3162]=8'b00110000;
    rom_data[3163]=rom_data[12];
    rom_data[3164]=8'b00110000;
    rom_data[3165]=rom_data[12];
    rom_data[3166]=8'b00110000;
    rom_data[3167]=rom_data[12];
    rom_data[3168]=8'b00110000;
    rom_data[3169]=rom_data[12];
    rom_data[3170]=8'b00110000;
    rom_data[3171]=rom_data[12];
    rom_data[3172]=8'b00110000;
    rom_data[3173]=rom_data[12];
    rom_data[3174]=8'b00110000;
    rom_data[3175]=rom_data[12];
    rom_data[3176]=8'b00110000;
    rom_data[3177]=rom_data[12];
    rom_data[3178]=8'b00110000;
    rom_data[3179]=rom_data[12];
    rom_data[3180]=8'b00101111;
    rom_data[3181]=rom_data[12];
    rom_data[3182]=8'b00101111;
    rom_data[3183]=rom_data[12];
    rom_data[3184]=8'b00101111;
    rom_data[3185]=rom_data[12];
    rom_data[3186]=8'b00101111;
    rom_data[3187]=rom_data[12];
    rom_data[3188]=8'b00101111;
    rom_data[3189]=rom_data[12];
    rom_data[3190]=8'b00101111;
    rom_data[3191]=rom_data[12];
    rom_data[3192]=8'b00101111;
    rom_data[3193]=rom_data[12];
    rom_data[3194]=8'b00101111;
    rom_data[3195]=rom_data[12];
    rom_data[3196]=8'b00101111;
    rom_data[3197]=rom_data[12];
    rom_data[3198]=8'b00101110;
    rom_data[3199]=rom_data[12];
    rom_data[3200]=8'b00101110;
    rom_data[3201]=rom_data[12];
    rom_data[3202]=8'b00101110;
    rom_data[3203]=rom_data[12];
    rom_data[3204]=8'b00101110;
    rom_data[3205]=rom_data[12];
    rom_data[3206]=8'b00101110;
    rom_data[3207]=rom_data[12];
    rom_data[3208]=8'b00101110;
    rom_data[3209]=rom_data[12];
    rom_data[3210]=8'b00101110;
    rom_data[3211]=rom_data[12];
    rom_data[3212]=8'b00101110;
    rom_data[3213]=rom_data[12];
    rom_data[3214]=8'b00101110;
    rom_data[3215]=rom_data[12];
    rom_data[3216]=8'b00101110;
    rom_data[3217]=rom_data[12];
    rom_data[3218]=8'b00101110;
    rom_data[3219]=rom_data[12];
    rom_data[3220]=8'b00101110;
    rom_data[3221]=rom_data[12];
    rom_data[3222]=8'b00101110;
    rom_data[3223]=rom_data[12];
    rom_data[3224]=8'b00101110;
    rom_data[3225]=rom_data[12];
    rom_data[3226]=8'b00101101;
    rom_data[3227]=rom_data[12];
    rom_data[3228]=8'b00101101;
    rom_data[3229]=rom_data[12];
    rom_data[3230]=8'b00101101;
    rom_data[3231]=rom_data[12];
    rom_data[3232]=8'b00101101;
    rom_data[3233]=rom_data[12];
    rom_data[3234]=8'b00101101;
    rom_data[3235]=rom_data[12];
    rom_data[3236]=8'b00101101;
    rom_data[3237]=rom_data[12];
    rom_data[3238]=8'b00101101;
    rom_data[3239]=rom_data[12];
    rom_data[3240]=8'b00101101;
    rom_data[3241]=rom_data[12];

  // F1   
  if (f1_addr==0) begin
    f1_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f1_addr==1) begin
    f1_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f1_addr[0]==1'b0) begin
    f1_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_D_q};
            end
            default: begin
            end
        endcase
   end // if addr=0
  // F2
  if (f2_addr==0) begin
    f2_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f2_addr==1) begin
    f2_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f2_addr[0]==1'b0) begin
    f2_data_d = 24'b00111000_0000000000000000; // Vref send in 50% samples  
  end else begin //data in 50%
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_D_q};
            end
            default: begin
            end
        endcase
   end // if addr=0
  // F3
  if (f3_addr==0) begin
    f3_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f3_addr==1) begin
    f3_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f3_addr[0]==1'b0) begin
    f3_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F4
  if (f4_addr==0) begin
    f4_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f4_addr==1) begin
    f4_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f4_addr[0]==1'b0) begin
    f4_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F5
  if (f5_addr==0) begin
    f5_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f5_addr==1) begin
    f5_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f5_addr[0]==1'b0) begin
    f5_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F6
  if (f6_addr==0) begin
    f6_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f6_addr==1) begin
    f6_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f6_addr[0]==1'b0) begin
    f6_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
end // always

always @(posedge f1_addr[0]) begin
    f1_CH_A_q<=f1_CH_A_d;
    f1_CH_B_q<=f1_CH_B_d;
    f1_CH_C_q<=f1_CH_C_d;
    f1_CH_D_q<=f1_CH_D_d;
end

always @(posedge f2_addr[0]) begin
    f2_CH_A_q<=f2_CH_A_d;
    f2_CH_B_q<=f2_CH_B_d;
    f2_CH_C_q<=f2_CH_C_d;
    f2_CH_D_q<=f2_CH_D_d;
end

always @(posedge f3_addr[0]) begin
    f3_CH_A_q<=f3_CH_A_d;
    f3_CH_B_q<=f3_CH_B_d;
    f3_CH_C_q<=f3_CH_C_d;
    f3_CH_D_q<=f3_CH_D_d;
end

always @(posedge f4_addr[0]) begin
    f4_CH_A_q<=f4_CH_A_d;
    f4_CH_B_q<=f4_CH_B_d;
    f4_CH_C_q<=f4_CH_C_d;
    f4_CH_D_q<=f4_CH_D_d;
end

always @(posedge f5_addr[0]) begin
    f5_CH_A_q<=f5_CH_A_d;
    f5_CH_B_q<=f5_CH_B_d;
    f5_CH_C_q<=f5_CH_C_d;
    f5_CH_D_q<=f5_CH_D_d;
end

always @(posedge f6_addr[0]) begin
    f6_CH_A_q<=f6_CH_A_d;
    f6_CH_B_q<=f6_CH_B_d;
    f6_CH_C_q<=f6_CH_C_d;
    f6_CH_D_q<=f6_CH_D_d;
end

always @(posedge clk) begin
    f1_data_q <= f1_data_d;
    f2_data_q <= f2_data_d;
    f3_data_q <= f3_data_d;
    f4_data_q <= f4_data_d;
    f5_data_q <= f5_data_d;
    f6_data_q <= f6_data_d;
end // always
 
endmodule