module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] f1_addr,
    input [15:0] f2_addr,
    input [15:0] f3_addr,
    input [15:0] f4_addr,
    input [15:0] f5_addr,
    input [15:0] f6_addr,

    input go_home,
    // OUTPUT
    output [23:0] f1_data,
    output [23:0] f2_data,
    output [23:0] f3_data,
    output [23:0] f4_data,
    output [23:0] f5_data,
    output [23:0] f6_data
    // output rom_scan_is_done
  );
  
parameter rom_size = 2201;

reg [15:0] rom_data [rom_size:0];

reg [23:0] f1_data_d, f1_data_q;
wire[13:0] f1_addrs;
reg [15:0] f1_antidata;

reg [23:0] f2_data_d, f2_data_q;
wire[13:0] f2_addrs;
reg [15:0] f2_antidata;

reg [23:0] f3_data_d, f3_data_q;
wire[13:0] f3_addrs;
reg [15:0] f3_antidata;

reg [23:0] f4_data_d, f4_data_q;
wire[13:0] f4_addrs;
reg [15:0] f4_antidata;

reg [23:0] f5_data_d, f5_data_q;
wire[13:0] f5_addrs;
reg [15:0] f5_antidata;

reg [23:0] f6_data_d, f6_data_q;
wire[13:0] f6_addrs;
reg [15:0] f6_antidata;

reg done;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;

reg [15:0] f1_CH_A_d, f1_CH_A_q;
reg [15:0] f1_CH_B_d, f1_CH_B_q;
reg [15:0] f1_CH_C_d, f1_CH_C_q;
reg [15:0] f1_CH_D_d, f1_CH_D_q;

reg [15:0] f2_CH_A_d, f2_CH_A_q;
reg [15:0] f2_CH_B_d, f2_CH_B_q;
reg [15:0] f2_CH_C_d, f2_CH_C_q;
reg [15:0] f2_CH_D_d, f2_CH_D_q;

reg [15:0] f3_CH_A_d, f3_CH_A_q;
reg [15:0] f3_CH_B_d, f3_CH_B_q;
reg [15:0] f3_CH_C_d, f3_CH_C_q;
reg [15:0] f3_CH_D_d, f3_CH_D_q;

reg [15:0] f4_CH_A_d, f4_CH_A_q;
reg [15:0] f4_CH_B_d, f4_CH_B_q;
reg [15:0] f4_CH_C_d, f4_CH_C_q;
reg [15:0] f4_CH_D_d, f4_CH_D_q;

reg [15:0] f5_CH_A_d, f5_CH_A_q;
reg [15:0] f5_CH_B_d, f5_CH_B_q;
reg [15:0] f5_CH_C_d, f5_CH_C_q;
reg [15:0] f5_CH_D_d, f5_CH_D_q;

reg [15:0] f6_CH_A_d, f6_CH_A_q;
reg [15:0] f6_CH_B_d, f6_CH_B_q;
reg [15:0] f6_CH_C_d, f6_CH_C_q;
reg [15:0] f6_CH_D_d, f6_CH_D_q;


assign f1_data = f1_data_q;
assign f2_data = f2_data_q;
assign f3_data = f3_data_q;
assign f4_data = f4_data_q;
assign f5_data = f5_data_q;
assign f6_data = f6_data_q;
// assign rom_scan_is_done = done;
assign f1_addrs = f1_addr[15:2];
assign f2_addrs = f2_addr[15:2];
assign f3_addrs = f3_addr[15:2];
assign f4_addrs = f4_addr[15:2];
assign f5_addrs = f5_addr[15:2];
assign f6_addrs = f6_addr[15:2];

always @(*) begin

    f1_CH_A_d=f1_CH_A_q;
    f1_CH_B_d=f1_CH_B_q;
    f1_CH_C_d=f1_CH_C_q;
    f1_CH_D_d=f1_CH_D_q;

    f2_CH_A_d=f2_CH_A_q;
    f2_CH_B_d=f2_CH_B_q;
    f2_CH_C_d=f2_CH_C_q;
    f2_CH_D_d=f2_CH_D_q;
    
    f3_CH_A_d=f3_CH_A_q;
    f3_CH_B_d=f3_CH_B_q;
    f3_CH_C_d=f3_CH_C_q;
    f3_CH_D_d=f3_CH_D_q;
    
    f4_CH_A_d=f4_CH_A_q;
    f4_CH_B_d=f4_CH_B_q;
    f4_CH_C_d=f4_CH_C_q;
    f4_CH_D_d=f4_CH_D_q;
    
    f5_CH_A_d=f5_CH_A_q;
    f5_CH_B_d=f5_CH_B_q;
    f5_CH_C_d=f5_CH_C_q;
    f5_CH_D_d=f5_CH_D_q;
    
    f6_CH_A_d=f6_CH_A_q;
    f6_CH_B_d=f6_CH_B_q;
    f6_CH_C_d=f6_CH_C_q;
    f6_CH_D_d=f6_CH_D_q;


    if (go_home==1'b1) begin
       
        // F1
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f1_CH_A_q>home_bias) begin
                    f1_CH_A_d=f1_CH_A_q-home_step;
                end else if (f1_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_A_d=f1_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f1_CH_C_q>home_bias) begin
                    f1_CH_C_d=f1_CH_C_q-home_step;
                end else if (f1_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_C_d=f1_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f1_CH_B_q>home_bias) begin
                    f1_CH_B_d=f1_CH_B_q-home_step;
                end else if (f1_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_B_d=f1_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f1_CH_D_q>home_bias) begin
                    f1_CH_D_d=f1_CH_D_q-home_step;
                end else if (f1_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_D_d=f1_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        
        // F2
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f2_CH_A_q>home_bias) begin
                    f2_CH_A_d=f2_CH_A_q-home_step;
                end else if (f2_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_A_d=f2_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f2_CH_C_q>home_bias) begin
                    f2_CH_C_d=f2_CH_C_q-home_step;
                end else if (f2_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_C_d=f2_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f2_CH_B_q>home_bias) begin
                    f2_CH_B_d=f2_CH_B_q-home_step;
                end else if (f2_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_B_d=f2_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f2_CH_D_q>home_bias) begin
                    f2_CH_D_d=f2_CH_D_q-home_step;
                end else if (f2_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_D_d=f2_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        
        // F3
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f3_CH_A_q>home_bias) begin
                    f3_CH_A_d=f3_CH_A_q-home_step;
                end else if (f3_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_A_d=f3_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f3_CH_C_q>home_bias) begin
                    f3_CH_C_d=f3_CH_C_q-home_step;
                end else if (f3_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_C_d=f3_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f3_CH_B_q>home_bias) begin
                    f3_CH_B_d=f3_CH_B_q-home_step;
                end else if (f3_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_B_d=f3_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f3_CH_D_q>home_bias) begin
                    f3_CH_D_d=f3_CH_D_q-home_step;
                end else if (f3_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_D_d=f3_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase

        // F4
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f4_CH_A_q>home_bias) begin
                    f4_CH_A_d=f4_CH_A_q-home_step;
                end else if (f4_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_A_d=f4_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f4_CH_C_q>home_bias) begin
                    f4_CH_C_d=f4_CH_C_q-home_step;
                end else if (f4_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_C_d=f4_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f4_CH_B_q>home_bias) begin
                    f4_CH_B_d=f4_CH_B_q-home_step;
                end else if (f4_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_B_d=f4_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f4_CH_D_q>home_bias) begin
                    f4_CH_D_d=f4_CH_D_q-home_step;
                end else if (f4_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_D_d=f4_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase

        // F5
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f5_CH_A_q>home_bias) begin
                    f5_CH_A_d=f5_CH_A_q-home_step;
                end else if (f5_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_A_d=f5_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f5_CH_C_q>home_bias) begin
                    f5_CH_C_d=f5_CH_C_q-home_step;
                end else if (f5_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_C_d=f5_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f5_CH_B_q>home_bias) begin
                    f5_CH_B_d=f5_CH_B_q-home_step;
                end else if (f5_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_B_d=f5_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f5_CH_D_q>home_bias) begin
                    f5_CH_D_d=f5_CH_D_q-home_step;
                end else if (f5_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_D_d=f5_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase

        // F6
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f6_CH_A_q>home_bias) begin
                    f6_CH_A_d=f6_CH_A_q-home_step;
                end else if (f6_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_A_d=f6_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f6_CH_C_q>home_bias) begin
                    f6_CH_C_d=f6_CH_C_q-home_step;
                end else if (f6_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_C_d=f6_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f6_CH_B_q>home_bias) begin
                    f6_CH_B_d=f6_CH_B_q-home_step;
                end else if (f6_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_B_d=f6_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f6_CH_D_q>home_bias) begin
                    f6_CH_D_d=f6_CH_D_q-home_step;
                end else if (f6_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_D_d=f6_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase

    end else begin // if go home==0
        
        // F1
        case (f1_addr[2:1])
            2'b00: begin
                f1_CH_A_d= rom_data[f1_addrs];
            end
            2'b01: begin
                f1_CH_C_d= f1_antidata;
            end
            2'b10: begin
                f1_CH_B_d= rom_data[f1_addrs];
            end
            2'b11: begin
                f1_CH_D_d= f1_antidata;
            end
        default: begin
            end
        endcase


        // F2
        case (f2_addr[2:1])
            2'b00: begin
                f2_CH_A_d= rom_data[f2_addrs];
            end
            2'b01: begin
                f2_CH_C_d= f2_antidata;
            end
            2'b10: begin
                f2_CH_B_d= rom_data[f2_addrs];
            end
            2'b11: begin
                f2_CH_D_d= f2_antidata;
            end
        default: begin
            end
        endcase

        // F3
        case (f3_addr[2:1])
            2'b00: begin
                f3_CH_A_d= rom_data[f3_addrs];
            end
            2'b01: begin
                f3_CH_C_d= f3_antidata;
            end
            2'b10: begin
                f3_CH_B_d= rom_data[f3_addrs];
            end
            2'b11: begin
                f3_CH_D_d= f3_antidata;
            end
        default: begin
            end
        endcase

        // F4
        case (f4_addr[2:1])
            2'b00: begin
                f4_CH_A_d= rom_data[f4_addrs];
            end
            2'b01: begin
                f4_CH_C_d= f4_antidata;
            end
            2'b10: begin
                f4_CH_B_d= rom_data[f4_addrs];
            end
            2'b11: begin
                f4_CH_D_d= f4_antidata;
            end
        default: begin
            end
        endcase

        // F5
        case (f5_addr[2:1])
            2'b00: begin
                f5_CH_A_d= rom_data[f5_addrs];
            end
            2'b01: begin
                f5_CH_C_d= f5_antidata;
            end
            2'b10: begin
                f5_CH_B_d= rom_data[f5_addrs];
            end
            2'b11: begin
                f5_CH_D_d= f5_antidata;
            end
        default: begin
            end
        endcase

        // F6
        case (f6_addr[2:1])
            2'b00: begin
                f6_CH_A_d= rom_data[f6_addrs];
            end
            2'b01: begin
                f6_CH_C_d= f6_antidata;
            end
            2'b10: begin
                f6_CH_B_d= rom_data[f6_addrs];
            end
            2'b11: begin
                f6_CH_D_d= f6_antidata;
            end
        default: begin
            end
        endcase


    end // if go home 



end // always





always @(*) begin
  f1_antidata = 16'hB900 - rom_data[f1_addrs];
  f2_antidata = 16'hB900 - rom_data[f2_addrs];
  f3_antidata = 16'hB900 - rom_data[f3_addrs];
  f4_antidata = 16'hB900 - rom_data[f4_addrs];
  f5_antidata = 16'hB900 - rom_data[f5_addrs];
  f6_antidata = 16'hB900 - rom_data[f6_addrs];
       
       
       

    rom_data[ 2]=16'b0011000001101101;
    rom_data[ 3]=16'b0101110111000000;
    rom_data[ 4]=16'b0011000010001000;
    rom_data[ 5]=16'b0101111011100111;
    rom_data[ 6]=16'b0011000010100011;
    rom_data[ 7]=16'b0110000000001101;
    rom_data[ 8]=16'b0011000010111111;
    rom_data[ 9]=16'b0110000100110011;
    rom_data[10]=16'b0011000011011011;
    rom_data[11]=16'b0110001001011001;
    rom_data[12]=16'b0011000011111001;
    rom_data[13]=16'b0110001101111111;
    rom_data[14]=16'b0011000100010111;
    rom_data[15]=16'b0110010010100100;
    rom_data[16]=16'b0011000100110110;
    rom_data[17]=16'b0110010111001001;
    rom_data[18]=16'b0011000101010101;
    rom_data[19]=16'b0110011011101100;
    rom_data[20]=16'b0011000101110101;
    rom_data[21]=16'b0110100000010000;
    rom_data[22]=16'b0011000110010110;
    rom_data[23]=16'b0110100100110010;
    rom_data[24]=16'b0011000110110111;
    rom_data[25]=16'b0110101001010011;
    rom_data[26]=16'b0011000111011001;
    rom_data[27]=16'b0110101101110011;
    rom_data[28]=16'b0011000111111011;
    rom_data[29]=16'b0110110010010010;
    rom_data[30]=16'b0011001000011110;
    rom_data[31]=16'b0110110110101111;
    rom_data[32]=16'b0011001001000001;
    rom_data[33]=16'b0110111011001100;
    rom_data[34]=16'b0011001001100101;
    rom_data[35]=16'b0110111111100110;
    rom_data[36]=16'b0011001010001010;
    rom_data[37]=16'b0111000011111111;
    rom_data[38]=16'b0011001010101110;
    rom_data[39]=16'b0111001000010110;
    rom_data[40]=16'b0011001011010100;
    rom_data[41]=16'b0111001100101100;
    rom_data[42]=16'b0011001011111010;
    rom_data[43]=16'b0111010000111111;
    rom_data[44]=16'b0011001100100000;
    rom_data[45]=16'b0111010101001111;
    rom_data[46]=16'b0011001101000111;
    rom_data[47]=16'b0111011001011110;
    rom_data[48]=16'b0011001101101111;
    rom_data[49]=16'b0111011101101010;
    rom_data[50]=16'b0011001110010110;
    rom_data[51]=16'b0111100001110011;
    rom_data[52]=16'b0011001110111111;
    rom_data[53]=16'b0111100101111001;
    rom_data[54]=16'b0011001111101000;
    rom_data[55]=16'b0111101001111100;
    rom_data[56]=16'b0011010000010010;
    rom_data[57]=16'b0111101101111100;
    rom_data[58]=16'b0011010000111100;
    rom_data[59]=16'b0111110001111000;
    rom_data[60]=16'b0011010001100110;
    rom_data[61]=16'b0111110101110000;
    rom_data[62]=16'b0011010010010010;
    rom_data[63]=16'b0111111001100100;
    rom_data[64]=16'b0011010010111101;
    rom_data[65]=16'b0111111101010011;
    rom_data[66]=16'b0011010011101010;
    rom_data[67]=16'b1000000000111110;
    rom_data[68]=16'b0011010100010111;
    rom_data[69]=16'b1000000100100100;
    rom_data[70]=16'b0011010101000100;
    rom_data[71]=16'b1000001000000101;
    rom_data[72]=16'b0011010101110011;
    rom_data[73]=16'b1000001011100000;
    rom_data[74]=16'b0011010110100001;
    rom_data[75]=16'b1000001110110101;
    rom_data[76]=16'b0011010111010001;
    rom_data[77]=16'b1000010010000011;
    rom_data[78]=16'b0011011000000001;
    rom_data[79]=16'b1000010101001011;
    rom_data[80]=16'b0011011000110001;
    rom_data[81]=16'b1000011000001100;
    rom_data[82]=16'b0011011001100010;
    rom_data[83]=16'b1000011011000100;
    rom_data[84]=16'b0011011010010100;
    rom_data[85]=16'b1000011101110101;
    rom_data[86]=16'b0011011011000110;
    rom_data[87]=16'b1000100000011100;
    rom_data[88]=16'b0011011011111001;
    rom_data[89]=16'b1000100010111011;
    rom_data[90]=16'b0011011100101100;
    rom_data[91]=16'b1000100101010000;
    rom_data[92]=16'b0011011101011111;
    rom_data[93]=16'b1000100111011010;
    rom_data[94]=16'b0011011110010011;
    rom_data[95]=16'b1000101001011010;
    rom_data[96]=16'b0011011111001000;
    rom_data[97]=16'b1000101011001110;
    rom_data[98]=16'b0011011111111100;
    rom_data[99]=16'b1000101100110110;
    rom_data[100]=16'b0011100000110001;
    rom_data[101]=16'b1000101110010010;
    rom_data[102]=16'b0011100001010101;
    rom_data[103]=16'b1000101111100001;
    rom_data[104]=16'b0011100010001011;
    rom_data[105]=16'b1000110000100011;
    rom_data[106]=16'b0011100011000000;
    rom_data[107]=16'b1000110001011000;
    rom_data[108]=16'b0011100011110110;
    rom_data[109]=16'b1000110001111110;
    rom_data[110]=16'b0011100100101100;
    rom_data[111]=16'b1000110010010110;
    rom_data[112]=16'b0011100101100001;
    rom_data[113]=16'b1000110010100000;
    rom_data[114]=16'b0011100110010110;
    rom_data[115]=16'b1000110010011011;
    rom_data[116]=16'b0011100111001010;
    rom_data[117]=16'b1000110010001000;
    rom_data[118]=16'b0011100111111111;
    rom_data[119]=16'b1000110001100110;
    rom_data[120]=16'b0011101000110011;
    rom_data[121]=16'b1000110000110111;
    rom_data[122]=16'b0011101001100110;
    rom_data[123]=16'b1000101111111001;
    rom_data[124]=16'b0011101010011001;
    rom_data[125]=16'b1000101110101110;
    rom_data[126]=16'b0011101011001100;
    rom_data[127]=16'b1000101101010101;
    rom_data[128]=16'b0011101011111110;
    rom_data[129]=16'b1000101011110000;
    rom_data[130]=16'b0011101100101111;
    rom_data[131]=16'b1000101001111110;
    rom_data[132]=16'b0011101101100000;
    rom_data[133]=16'b1000101000000001;
    rom_data[134]=16'b0011101110010001;
    rom_data[135]=16'b1000100101111000;
    rom_data[136]=16'b0011101111000001;
    rom_data[137]=16'b1000100011100101;
    rom_data[138]=16'b0011101111110000;
    rom_data[139]=16'b1000100001000111;
    rom_data[140]=16'b0011110000011111;
    rom_data[141]=16'b1000011110100000;
    rom_data[142]=16'b0011110001001110;
    rom_data[143]=16'b1000011011110000;
    rom_data[144]=16'b0011110001111100;
    rom_data[145]=16'b1000011000110111;
    rom_data[146]=16'b0011110010101001;
    rom_data[147]=16'b1000010101110110;
    rom_data[148]=16'b0011110011010110;
    rom_data[149]=16'b1000010010101110;
    rom_data[150]=16'b0011110100000011;
    rom_data[151]=16'b1000001111011111;
    rom_data[152]=16'b0011110100101111;
    rom_data[153]=16'b1000001100001001;
    rom_data[154]=16'b0011110101011010;
    rom_data[155]=16'b1000001000101101;
    rom_data[156]=16'b0011110110000110;
    rom_data[157]=16'b1000000101001011;
    rom_data[158]=16'b0011110110110001;
    rom_data[159]=16'b1000000001100011;
    rom_data[160]=16'b0011110111011011;
    rom_data[161]=16'b0111111101110111;
    rom_data[162]=16'b0011111000000101;
    rom_data[163]=16'b0111111010000101;
    rom_data[164]=16'b0011111000101111;
    rom_data[165]=16'b0111110110010000;
    rom_data[166]=16'b0011111001011001;
    rom_data[167]=16'b0111110010010110;
    rom_data[168]=16'b0011111010000010;
    rom_data[169]=16'b0111101110011000;
    rom_data[170]=16'b0011111010101011;
    rom_data[171]=16'b0111101010010111;
    rom_data[172]=16'b0011111011010100;
    rom_data[173]=16'b0111100110010010;
    rom_data[174]=16'b0011111011111100;
    rom_data[175]=16'b0111100010001010;
    rom_data[176]=16'b0011111100100100;
    rom_data[177]=16'b0111011101111111;
    rom_data[178]=16'b0011111101001100;
    rom_data[179]=16'b0111011001110010;
    rom_data[180]=16'b0011111101110100;
    rom_data[181]=16'b0111010101100010;
    rom_data[182]=16'b0011111110011011;
    rom_data[183]=16'b0111010001001111;
    rom_data[184]=16'b0011111111000011;
    rom_data[185]=16'b0111001100111011;
    rom_data[186]=16'b0011111111101010;
    rom_data[187]=16'b0111001000100100;
    rom_data[188]=16'b0100000000010001;
    rom_data[189]=16'b0111000100001011;
    rom_data[190]=16'b0100000000111000;
    rom_data[191]=16'b0110111111110001;
    rom_data[192]=16'b0100000001011110;
    rom_data[193]=16'b0110111011010101;
    rom_data[194]=16'b0100000010000101;
    rom_data[195]=16'b0110110110111000;
    rom_data[196]=16'b0100000010101011;
    rom_data[197]=16'b0110110010011001;
    rom_data[198]=16'b0100000011010010;
    rom_data[199]=16'b0110101101111001;
    rom_data[200]=16'b0100000011111000;
    rom_data[201]=16'b0110101001011000;
    rom_data[202]=16'b0100000100011110;
    rom_data[203]=16'b0110100100110110;
    rom_data[204]=16'b0100000101000100;
    rom_data[205]=16'b0110100000010011;
    rom_data[206]=16'b0100000101101011;
    rom_data[207]=16'b0110011011101111;
    rom_data[208]=16'b0100000110010001;
    rom_data[209]=16'b0110010111001011;
    rom_data[210]=16'b0100000110110111;
    rom_data[211]=16'b0110010010100110;
    rom_data[212]=16'b0100000111011101;
    rom_data[213]=16'b0110001110000000;
    rom_data[214]=16'b0100001000000011;
    rom_data[215]=16'b0110001001011010;
    rom_data[216]=16'b0100001000101001;
    rom_data[217]=16'b0110000100110100;
    rom_data[218]=16'b0100001001001111;
    rom_data[219]=16'b0110000000001101;
    rom_data[220]=16'b0100001001110101;
    rom_data[221]=16'b0101111011100111;
    rom_data[222]=16'b0100001010011011;
    rom_data[223]=16'b0101110111000000;
    rom_data[224]=16'b0100001011000001;
    rom_data[225]=16'b0101110010011001;
    rom_data[226]=16'b0100001011100111;
    rom_data[227]=16'b0101101101110011;
    rom_data[228]=16'b0100001100001101;
    rom_data[229]=16'b0101101001001100;
    rom_data[230]=16'b0100001100110100;
    rom_data[231]=16'b0101100100100110;
    rom_data[232]=16'b0100001101011010;
    rom_data[233]=16'b0101100000000001;
    rom_data[234]=16'b0100001110000001;
    rom_data[235]=16'b0101011011011100;
    rom_data[236]=16'b0100001110100111;
    rom_data[237]=16'b0101010110110111;
    rom_data[238]=16'b0100001111001110;
    rom_data[239]=16'b0101010010010011;
    rom_data[240]=16'b0100001111110101;
    rom_data[241]=16'b0101001101110000;
    rom_data[242]=16'b0100010000011100;
    rom_data[243]=16'b0101001001001110;
    rom_data[244]=16'b0100010001000100;
    rom_data[245]=16'b0101000100101101;
    rom_data[246]=16'b0100010001101011;
    rom_data[247]=16'b0101000000001101;
    rom_data[248]=16'b0100010010010011;
    rom_data[249]=16'b0100111011101110;
    rom_data[250]=16'b0100010010111011;
    rom_data[251]=16'b0100110111010000;
    rom_data[252]=16'b0100010011100011;
    rom_data[253]=16'b0100110010110100;
    rom_data[254]=16'b0100010100001011;
    rom_data[255]=16'b0100101110011010;
    rom_data[256]=16'b0100010100110100;
    rom_data[257]=16'b0100101010000001;
    rom_data[258]=16'b0100010101011101;
    rom_data[259]=16'b0100100101101010;
    rom_data[260]=16'b0100010110000110;
    rom_data[261]=16'b0100100001010100;
    rom_data[262]=16'b0100010110110000;
    rom_data[263]=16'b0100011101000001;
    rom_data[264]=16'b0100010111011001;
    rom_data[265]=16'b0100011000110000;
    rom_data[266]=16'b0100011000000100;
    rom_data[267]=16'b0100010100100010;
    rom_data[268]=16'b0100011000101110;
    rom_data[269]=16'b0100010000010110;
    rom_data[270]=16'b0100011001011001;
    rom_data[271]=16'b0100001100001101;
    rom_data[272]=16'b0100011010000100;
    rom_data[273]=16'b0100001000000111;
    rom_data[274]=16'b0100011010110000;
    rom_data[275]=16'b0100000100000100;
    rom_data[276]=16'b0100011011011100;
    rom_data[277]=16'b0100000000000100;
    rom_data[278]=16'b0100011100001000;
    rom_data[279]=16'b0011111100001000;
    rom_data[280]=16'b0100011100110101;
    rom_data[281]=16'b0011111000010000;
    rom_data[282]=16'b0100011101100011;
    rom_data[283]=16'b0011110100011100;
    rom_data[284]=16'b0100011110010001;
    rom_data[285]=16'b0011110000101100;
    rom_data[286]=16'b0100011110111111;
    rom_data[287]=16'b0011101101000010;
    rom_data[288]=16'b0100011111101110;
    rom_data[289]=16'b0011101001011100;
    rom_data[290]=16'b0100100000011101;
    rom_data[291]=16'b0011100101111011;
    rom_data[292]=16'b0100100001001101;
    rom_data[293]=16'b0011100010100000;
    rom_data[294]=16'b0100100001111101;
    rom_data[295]=16'b0011011111001011;
    rom_data[296]=16'b0100100010101110;
    rom_data[297]=16'b0011011011111100;
    rom_data[298]=16'b0100100011100000;
    rom_data[299]=16'b0011011000110101;
    rom_data[300]=16'b0100100100010010;
    rom_data[301]=16'b0011010101110100;
    rom_data[302]=16'b0100100101000100;
    rom_data[303]=16'b0011010010111100;
    rom_data[304]=16'b0100100101110111;
    rom_data[305]=16'b0011010000001011;
    rom_data[306]=16'b0100100110101010;
    rom_data[307]=16'b0011001101100100;
    rom_data[308]=16'b0100100111011110;
    rom_data[309]=16'b0011001011000101;
    rom_data[310]=16'b0100101000010010;
    rom_data[311]=16'b0011001000110000;
    rom_data[312]=16'b0100101001000111;
    rom_data[313]=16'b0011000110100110;
    rom_data[314]=16'b0100101001111100;
    rom_data[315]=16'b0011000100100110;
    rom_data[316]=16'b0100101010110001;
    rom_data[317]=16'b0011000010110010;
    rom_data[318]=16'b0100101011100110;
    rom_data[319]=16'b0011000001001010;
    rom_data[320]=16'b0100101100011100;
    rom_data[321]=16'b0010111111101110;
    rom_data[322]=16'b0100101101010010;
    rom_data[323]=16'b0010111110011110;
    rom_data[324]=16'b0100101110000111;
    rom_data[325]=16'b0010111101011101;
    rom_data[326]=16'b0100101110111101;
    rom_data[327]=16'b0010111100101000;
    rom_data[328]=16'b0100101111110011;
    rom_data[329]=16'b0010111100000010;
    rom_data[330]=16'b0100110000101000;
    rom_data[331]=16'b0010111011101010;
    rom_data[332]=16'b0100110001011101;
    rom_data[333]=16'b0010111011100000;
    rom_data[334]=16'b0100110010010010;
    rom_data[335]=16'b0010111011100101;
    rom_data[336]=16'b0100110011000111;
    rom_data[337]=16'b0010111011111000;
    rom_data[338]=16'b0100110011111011;
    rom_data[339]=16'b0010111100011010;
    rom_data[340]=16'b0100110100101111;
    rom_data[341]=16'b0010111101001001;
    rom_data[342]=16'b0100110101100011;
    rom_data[343]=16'b0010111110000111;
    rom_data[344]=16'b0100110110010110;
    rom_data[345]=16'b0010111111010010;
    rom_data[346]=16'b0100110111001000;
    rom_data[347]=16'b0011000000101011;
    rom_data[348]=16'b0100110111111010;
    rom_data[349]=16'b0011000010010000;
    rom_data[350]=16'b0100111000101100;
    rom_data[351]=16'b0011000100000010;
    rom_data[352]=16'b0100111001011101;
    rom_data[353]=16'b0011000101111111;
    rom_data[354]=16'b0100111010001101;
    rom_data[355]=16'b0011001000001000;
    rom_data[356]=16'b0100111010111101;
    rom_data[357]=16'b0011001010011011;
    rom_data[358]=16'b0100111011101101;
    rom_data[359]=16'b0011001100111001;
    rom_data[360]=16'b0100111100011100;
    rom_data[361]=16'b0011001111100000;
    rom_data[362]=16'b0100111101001010;
    rom_data[363]=16'b0011010010010000;
    rom_data[364]=16'b0100111101111000;
    rom_data[365]=16'b0011010101001001;
    rom_data[366]=16'b0100111110100110;
    rom_data[367]=16'b0011011000001010;
    rom_data[368]=16'b0100111111010011;
    rom_data[369]=16'b0011011011010010;
    rom_data[370]=16'b0100111111111111;
    rom_data[371]=16'b0011011110100001;
    rom_data[372]=16'b0101000000101011;
    rom_data[373]=16'b0011100001110111;
    rom_data[374]=16'b0101000001010111;
    rom_data[375]=16'b0011100101010011;
    rom_data[376]=16'b0101000010000010;
    rom_data[377]=16'b0011101000110101;
    rom_data[378]=16'b0101000010101101;
    rom_data[379]=16'b0011101100011101;
    rom_data[380]=16'b0101000011011000;
    rom_data[381]=16'b0011110000001001;
    rom_data[382]=16'b0101000100000010;
    rom_data[383]=16'b0011110011111011;
    rom_data[384]=16'b0101000100101100;
    rom_data[385]=16'b0011110111110000;
    rom_data[386]=16'b0101000101010101;
    rom_data[387]=16'b0011111011101010;
    rom_data[388]=16'b0101000101111111;
    rom_data[389]=16'b0011111111101000;
    rom_data[390]=16'b0101000110101000;
    rom_data[391]=16'b0100000011101001;
    rom_data[392]=16'b0101000111010000;
    rom_data[393]=16'b0100000111101110;
    rom_data[394]=16'b0101000111111001;
    rom_data[395]=16'b0100001011110110;
    rom_data[396]=16'b0101001000100001;
    rom_data[397]=16'b0100010000000001;
    rom_data[398]=16'b0101001001001001;
    rom_data[399]=16'b0100010100001110;
    rom_data[400]=16'b0101001001110000;
    rom_data[401]=16'b0100011000011110;
    rom_data[402]=16'b0101001010011000;
    rom_data[403]=16'b0100011100110001;
    rom_data[404]=16'b0101001010111111;
    rom_data[405]=16'b0100100001000101;
    rom_data[406]=16'b0101001011100110;
    rom_data[407]=16'b0100100101011100;
    rom_data[408]=16'b0101001100001101;
    rom_data[409]=16'b0100101001110101;
    rom_data[410]=16'b0101001100110100;
    rom_data[411]=16'b0100101110001111;
    rom_data[412]=16'b0101001101011011;
    rom_data[413]=16'b0100110010101011;
    rom_data[414]=16'b0101001110000010;
    rom_data[415]=16'b0100110111001000;
    rom_data[416]=16'b0101001110101000;
    rom_data[417]=16'b0100111011100111;
    rom_data[418]=16'b0101001111001110;
    rom_data[419]=16'b0101000000000111;
    rom_data[420]=16'b0101001111110101;
    rom_data[421]=16'b0101000100101000;
    rom_data[422]=16'b0101010000011011;
    rom_data[423]=16'b0101001001001010;
    rom_data[424]=16'b0101010001000001;
    rom_data[425]=16'b0101001101101101;
    rom_data[426]=16'b0101010001100111;
    rom_data[427]=16'b0101010010010001;
    rom_data[428]=16'b0101010010001101;
    rom_data[429]=16'b0101010110110101;
    rom_data[430]=16'b0101010010110011;
    rom_data[431]=16'b0101011011011011;
    rom_data[432]=16'b0101010011011001;
    rom_data[433]=16'b0101100000000000;
    rom_data[434]=16'b0101010011111111;
    rom_data[435]=16'b0101100100100110;
    rom_data[436]=16'b0101010100100101;
    rom_data[437]=16'b0101101001001100;
    rom_data[438]=16'b0101010101001011;
    rom_data[439]=16'b0101101101110011;
    rom_data[440]=16'b0101010101110001;
    rom_data[441]=16'b0101110010011010;
    rom_data[442]=16'b0101010110010111;
    rom_data[443]=16'b0101110111000000;
    rom_data[444]=16'b0101010110111101;
    rom_data[445]=16'b0101111011100111;
    rom_data[446]=16'b0101010111100100;
    rom_data[447]=16'b0110000000001101;
    rom_data[448]=16'b0101011000001010;
    rom_data[449]=16'b0110000100110100;
    rom_data[450]=16'b0101011000110000;
    rom_data[451]=16'b0110001001011010;
    rom_data[452]=16'b0101011001010111;
    rom_data[453]=16'b0110001101111111;
    rom_data[454]=16'b0101011001111101;
    rom_data[455]=16'b0110010010100100;
    rom_data[456]=16'b0101011010100100;
    rom_data[457]=16'b0110010111001001;
    rom_data[458]=16'b0101011011001011;
    rom_data[459]=16'b0110011011101101;
    rom_data[460]=16'b0101011011110010;
    rom_data[461]=16'b0110100000010000;
    rom_data[462]=16'b0101011100011001;
    rom_data[463]=16'b0110100100110010;
    rom_data[464]=16'b0101011101000000;
    rom_data[465]=16'b0110101001010011;
    rom_data[466]=16'b0101011101101000;
    rom_data[467]=16'b0110101101110011;
    rom_data[468]=16'b0101011110001111;
    rom_data[469]=16'b0110110010010010;
    rom_data[470]=16'b0101011110110111;
    rom_data[471]=16'b0110110110110000;
    rom_data[472]=16'b0101011111100000;
    rom_data[473]=16'b0110111011001100;
    rom_data[474]=16'b0101100000001000;
    rom_data[475]=16'b0110111111100111;
    rom_data[476]=16'b0101100000110001;
    rom_data[477]=16'b0111000100000000;
    rom_data[478]=16'b0101100001011001;
    rom_data[479]=16'b0111001000010111;
    rom_data[480]=16'b0101100010000011;
    rom_data[481]=16'b0111001100101100;
    rom_data[482]=16'b0101100010101100;
    rom_data[483]=16'b0111010000111111;
    rom_data[484]=16'b0101100011010110;
    rom_data[485]=16'b0111010101010000;
    rom_data[486]=16'b0101100100000000;
    rom_data[487]=16'b0111011001011110;
    rom_data[488]=16'b0101100100101011;
    rom_data[489]=16'b0111011101101010;
    rom_data[490]=16'b0101100101010110;
    rom_data[491]=16'b0111100001110011;
    rom_data[492]=16'b0101100110000001;
    rom_data[493]=16'b0111100101111001;
    rom_data[494]=16'b0101100110101100;
    rom_data[495]=16'b0111101001111100;
    rom_data[496]=16'b0101100111011001;
    rom_data[497]=16'b0111101101111100;
    rom_data[498]=16'b0101101000000101;
    rom_data[499]=16'b0111110001111000;
    rom_data[500]=16'b0101101000110010;
    rom_data[501]=16'b0111110101110000;
    rom_data[502]=16'b0101101001011111;
    rom_data[503]=16'b0111111001100100;
    rom_data[504]=16'b0101101010001101;
    rom_data[505]=16'b0111111101010100;
    rom_data[506]=16'b0101101010111100;
    rom_data[507]=16'b1000000000111111;
    rom_data[508]=16'b0101101011101010;
    rom_data[509]=16'b1000000100100101;
    rom_data[510]=16'b0101101100011010;
    rom_data[511]=16'b1000001000000101;
    rom_data[512]=16'b0101101101001010;
    rom_data[513]=16'b1000001011100000;
    rom_data[514]=16'b0101101101111010;
    rom_data[515]=16'b1000001110110101;
    rom_data[516]=16'b0101101110101011;
    rom_data[517]=16'b1000010010000100;
    rom_data[518]=16'b0101101111011100;
    rom_data[519]=16'b1000010101001011;
    rom_data[520]=16'b0101110000001110;
    rom_data[521]=16'b1000011000001100;
    rom_data[522]=16'b0101110001000001;
    rom_data[523]=16'b1000011011000100;
    rom_data[524]=16'b0101110001110011;
    rom_data[525]=16'b1000011101110101;
    rom_data[526]=16'b0101110010100111;
    rom_data[527]=16'b1000100000011101;
    rom_data[528]=16'b0101110011011011;
    rom_data[529]=16'b1000100010111011;
    rom_data[530]=16'b0101110100001111;
    rom_data[531]=16'b1000100101010000;
    rom_data[532]=16'b0101110101000011;
    rom_data[533]=16'b1000100111011010;
    rom_data[534]=16'b0101110101111000;
    rom_data[535]=16'b1000101001011010;
    rom_data[536]=16'b0101110110101101;
    rom_data[537]=16'b1000101011001110;
    rom_data[538]=16'b0101110111100011;
    rom_data[539]=16'b1000101100110110;
    rom_data[540]=16'b0101111000011000;
    rom_data[541]=16'b1000101110010010;
    rom_data[542]=16'b0101111001001110;
    rom_data[543]=16'b1000101111100010;
    rom_data[544]=16'b0101111010000100;
    rom_data[545]=16'b1000110000100011;
    rom_data[546]=16'b0101111010111010;
    rom_data[547]=16'b1000110001011000;
    rom_data[548]=16'b0101111011101111;
    rom_data[549]=16'b1000110001111110;
    rom_data[550]=16'b0101111100100101;
    rom_data[551]=16'b1000110010010110;
    rom_data[552]=16'b0101111101011010;
    rom_data[553]=16'b1000110010100000;
    rom_data[554]=16'b0101111110001111;
    rom_data[555]=16'b1000110010011011;
    rom_data[556]=16'b0101111111000100;
    rom_data[557]=16'b1000110010001000;
    rom_data[558]=16'b0101111111111000;
    rom_data[559]=16'b1000110001100110;
    rom_data[560]=16'b0110000000101100;
    rom_data[561]=16'b1000110000110111;
    rom_data[562]=16'b0110000001011111;
    rom_data[563]=16'b1000101111111001;
    rom_data[564]=16'b0110000010010010;
    rom_data[565]=16'b1000101110101101;
    rom_data[566]=16'b0110000011000101;
    rom_data[567]=16'b1000101101010101;
    rom_data[568]=16'b0110000011110111;
    rom_data[569]=16'b1000101011110000;
    rom_data[570]=16'b0110000100101001;
    rom_data[571]=16'b1000101001111110;
    rom_data[572]=16'b0110000101011010;
    rom_data[573]=16'b1000101000000001;
    rom_data[574]=16'b0110000110001010;
    rom_data[575]=16'b1000100101111000;
    rom_data[576]=16'b0110000110111010;
    rom_data[577]=16'b1000100011100101;
    rom_data[578]=16'b0110000111101001;
    rom_data[579]=16'b1000100001000111;
    rom_data[580]=16'b0110001000011000;
    rom_data[581]=16'b1000011110100000;
    rom_data[582]=16'b0110001001000111;
    rom_data[583]=16'b1000011011110000;
    rom_data[584]=16'b0110001001110101;
    rom_data[585]=16'b1000011000110111;
    rom_data[586]=16'b0110001010100010;
    rom_data[587]=16'b1000010101110110;
    rom_data[588]=16'b0110001011001111;
    rom_data[589]=16'b1000010010101110;
    rom_data[590]=16'b0110001011111100;
    rom_data[591]=16'b1000001111011111;
    rom_data[592]=16'b0110001100101000;
    rom_data[593]=16'b1000001100001001;
    rom_data[594]=16'b0110001101010100;
    rom_data[595]=16'b1000001000101100;
    rom_data[596]=16'b0110001101111111;
    rom_data[597]=16'b1000000101001010;
    rom_data[598]=16'b0110001110101010;
    rom_data[599]=16'b1000000001100011;
    rom_data[600]=16'b0110001111010100;
    rom_data[601]=16'b0111111101110110;
    rom_data[602]=16'b0110001111111111;
    rom_data[603]=16'b0111111010000101;
    rom_data[604]=16'b0110010000101000;
    rom_data[605]=16'b0111110110001111;
    rom_data[606]=16'b0110010001010010;
    rom_data[607]=16'b0111110010010110;
    rom_data[608]=16'b0110010001111011;
    rom_data[609]=16'b0111101110011000;
    rom_data[610]=16'b0110010010100100;
    rom_data[611]=16'b0111101010010111;
    rom_data[612]=16'b0110010011001101;
    rom_data[613]=16'b0111100110010010;
    rom_data[614]=16'b0110010011110101;
    rom_data[615]=16'b0111100010001010;
    rom_data[616]=16'b0110010100011101;
    rom_data[617]=16'b0111011101111111;
    rom_data[618]=16'b0110010101000101;
    rom_data[619]=16'b0111011001110010;
    rom_data[620]=16'b0110010101101101;
    rom_data[621]=16'b0111010101100010;
    rom_data[622]=16'b0110010110010101;
    rom_data[623]=16'b0111010001001111;
    rom_data[624]=16'b0110010110111100;
    rom_data[625]=16'b0111001100111010;
    rom_data[626]=16'b0110010111100011;
    rom_data[627]=16'b0111001000100100;
    rom_data[628]=16'b0110011000001010;
    rom_data[629]=16'b0111000100001011;
    rom_data[630]=16'b0110011000110001;
    rom_data[631]=16'b0110111111110001;
    rom_data[632]=16'b0110011001011000;
    rom_data[633]=16'b0110111011010101;
    rom_data[634]=16'b0110011001111110;
    rom_data[635]=16'b0110110110111000;
    rom_data[636]=16'b0110011010100101;
    rom_data[637]=16'b0110110010011001;
    rom_data[638]=16'b0110011011001011;
    rom_data[639]=16'b0110101101111001;
    rom_data[640]=16'b0110011011110001;
    rom_data[641]=16'b0110101001011000;
    rom_data[642]=16'b0110011100010111;
    rom_data[643]=16'b0110100100110110;
    rom_data[644]=16'b0110011100111110;
    rom_data[645]=16'b0110100000010011;
    rom_data[646]=16'b0110011101100100;
    rom_data[647]=16'b0110011011101111;
    rom_data[648]=16'b0110011110001010;
    rom_data[649]=16'b0110010111001010;
    rom_data[650]=16'b0110011110110000;
    rom_data[651]=16'b0110010010100101;
    rom_data[652]=16'b0110011111010110;
    rom_data[653]=16'b0110001110000000;
    rom_data[654]=16'b0110011111111100;
    rom_data[655]=16'b0110001001011010;
    rom_data[656]=16'b0110100000100010;
    rom_data[657]=16'b0110000100110011;
    rom_data[658]=16'b0110100001001000;
    rom_data[659]=16'b0110000000001101;
    rom_data[660]=16'b0110100001101110;
    rom_data[661]=16'b0101111011100110;
    rom_data[662]=16'b0110100010010100;
    rom_data[663]=16'b0101110111000000;
    rom_data[664]=16'b0110100010111010;
    rom_data[665]=16'b0101110010011001;
    rom_data[666]=16'b0110100011100000;
    rom_data[667]=16'b0101101101110010;
    rom_data[668]=16'b0110100100000110;
    rom_data[669]=16'b0101101001001100;
    rom_data[670]=16'b0110100100101101;
    rom_data[671]=16'b0101100100100110;
    rom_data[672]=16'b0110100101010011;
    rom_data[673]=16'b0101100000000000;
    rom_data[674]=16'b0110100101111010;
    rom_data[675]=16'b0101011011011011;
    rom_data[676]=16'b0110100110100001;
    rom_data[677]=16'b0101010110110111;
    rom_data[678]=16'b0110100111000111;
    rom_data[679]=16'b0101010010010011;
    rom_data[680]=16'b0110100111101110;
    rom_data[681]=16'b0101001101110000;
    rom_data[682]=16'b0110101000010110;
    rom_data[683]=16'b0101001001001110;
    rom_data[684]=16'b0110101000111101;
    rom_data[685]=16'b0101000100101101;
    rom_data[686]=16'b0110101001100100;
    rom_data[687]=16'b0101000000001101;
    rom_data[688]=16'b0110101010001100;
    rom_data[689]=16'b0100111011101110;
    rom_data[690]=16'b0110101010110100;
    rom_data[691]=16'b0100110111010000;
    rom_data[692]=16'b0110101011011100;
    rom_data[693]=16'b0100110010110100;
    rom_data[694]=16'b0110101100000100;
    rom_data[695]=16'b0100101110011001;
    rom_data[696]=16'b0110101100101101;
    rom_data[697]=16'b0100101010000000;
    rom_data[698]=16'b0110101101010110;
    rom_data[699]=16'b0100100101101001;
    rom_data[700]=16'b0110101101111111;
    rom_data[701]=16'b0100100001010100;
    rom_data[702]=16'b0110101110101001;
    rom_data[703]=16'b0100011101000001;
    rom_data[704]=16'b0110101111010011;
    rom_data[705]=16'b0100011000110000;
    rom_data[706]=16'b0110101111111101;
    rom_data[707]=16'b0100010100100010;
    rom_data[708]=16'b0110110000100111;
    rom_data[709]=16'b0100010000010110;
    rom_data[710]=16'b0110110001010010;
    rom_data[711]=16'b0100001100001101;
    rom_data[712]=16'b0110110001111101;
    rom_data[713]=16'b0100001000000111;
    rom_data[714]=16'b0110110010101001;
    rom_data[715]=16'b0100000100000100;
    rom_data[716]=16'b0110110011010101;
    rom_data[717]=16'b0100000000000100;
    rom_data[718]=16'b0110110100000010;
    rom_data[719]=16'b0011111100001000;
    rom_data[720]=16'b0110110100101111;
    rom_data[721]=16'b0011111000010000;
    rom_data[722]=16'b0110110101011100;
    rom_data[723]=16'b0011110100011100;
    rom_data[724]=16'b0110110110001010;
    rom_data[725]=16'b0011110000101100;
    rom_data[726]=16'b0110110110111000;
    rom_data[727]=16'b0011101101000001;
    rom_data[728]=16'b0110110111100111;
    rom_data[729]=16'b0011101001011011;
    rom_data[730]=16'b0110111000010110;
    rom_data[731]=16'b0011100101111011;
    rom_data[732]=16'b0110111001000110;
    rom_data[733]=16'b0011100010100000;
    rom_data[734]=16'b0110111001110111;
    rom_data[735]=16'b0011011111001011;
    rom_data[736]=16'b0110111010100111;
    rom_data[737]=16'b0011011011111100;
    rom_data[738]=16'b0110111011011001;
    rom_data[739]=16'b0011011000110101;
    rom_data[740]=16'b0110111100001011;
    rom_data[741]=16'b0011010101110100;
    rom_data[742]=16'b0110111100111101;
    rom_data[743]=16'b0011010010111100;
    rom_data[744]=16'b0110111101110000;
    rom_data[745]=16'b0011010000001011;
    rom_data[746]=16'b0110111110100011;
    rom_data[747]=16'b0011001101100011;
    rom_data[748]=16'b0110111111010111;
    rom_data[749]=16'b0011001011000101;
    rom_data[750]=16'b0111000000001011;
    rom_data[751]=16'b0011001000110000;
    rom_data[752]=16'b0111000001000000;
    rom_data[753]=16'b0011000110100110;
    rom_data[754]=16'b0111000001110101;
    rom_data[755]=16'b0011000100100110;
    rom_data[756]=16'b0111000010101010;
    rom_data[757]=16'b0011000010110010;
    rom_data[758]=16'b0111000011011111;
    rom_data[759]=16'b0011000001001010;
    rom_data[760]=16'b0111000100010101;
    rom_data[761]=16'b0010111111101110;
    rom_data[762]=16'b0111000101001011;
    rom_data[763]=16'b0010111110011110;
    rom_data[764]=16'b0111000110000000;
    rom_data[765]=16'b0010111101011101;
    rom_data[766]=16'b0111000110110110;
    rom_data[767]=16'b0010111100101000;
    rom_data[768]=16'b0111000111101100;
    rom_data[769]=16'b0010111100000010;
    rom_data[770]=16'b0111001000100001;
    rom_data[771]=16'b0010111011101010;
    rom_data[772]=16'b0111001001010111;
    rom_data[773]=16'b0010111011100000;
    rom_data[774]=16'b0111001010001100;
    rom_data[775]=16'b0010111011100101;
    rom_data[776]=16'b0111001011000000;
    rom_data[777]=16'b0010111011111000;
    rom_data[778]=16'b0111001011110101;
    rom_data[779]=16'b0010111100011010;
    rom_data[780]=16'b0111001100101000;
    rom_data[781]=16'b0010111101001010;
    rom_data[782]=16'b0111001101011100;
    rom_data[783]=16'b0010111110000111;
    rom_data[784]=16'b0111001110001111;
    rom_data[785]=16'b0010111111010011;
    rom_data[786]=16'b0111001111000010;
    rom_data[787]=16'b0011000000101011;
    rom_data[788]=16'b0111001111110100;
    rom_data[789]=16'b0011000010010000;
    rom_data[790]=16'b0111010000100101;
    rom_data[791]=16'b0011000100000010;
    rom_data[792]=16'b0111010001010110;
    rom_data[793]=16'b0011000101111111;
    rom_data[794]=16'b0111010010000111;
    rom_data[795]=16'b0011001000001000;
    rom_data[796]=16'b0111010010110111;
    rom_data[797]=16'b0011001010011100;
    rom_data[798]=16'b0111010011100110;
    rom_data[799]=16'b0011001100111001;
    rom_data[800]=16'b0111010100010101;
    rom_data[801]=16'b0011001111100000;
    rom_data[802]=16'b0111010101000011;
    rom_data[803]=16'b0011010010010000;
    rom_data[804]=16'b0111010101110001;
    rom_data[805]=16'b0011010101001001;
    rom_data[806]=16'b0111010110011111;
    rom_data[807]=16'b0011011000001010;
    rom_data[808]=16'b0111010111001100;
    rom_data[809]=16'b0011011011010010;
    rom_data[810]=16'b0111010111111000;
    rom_data[811]=16'b0011011110100010;
    rom_data[812]=16'b0111011000100100;
    rom_data[813]=16'b0011100001110111;
    rom_data[814]=16'b0111011001010000;
    rom_data[815]=16'b0011100101010100;
    rom_data[816]=16'b0111011001111100;
    rom_data[817]=16'b0011101000110110;
    rom_data[818]=16'b0111011010100110;
    rom_data[819]=16'b0011101100011101;
    rom_data[820]=16'b0111011011010001;
    rom_data[821]=16'b0011110000001010;
    rom_data[822]=16'b0111011011111011;
    rom_data[823]=16'b0011110011111011;
    rom_data[824]=16'b0111011100100101;
    rom_data[825]=16'b0011110111110001;
    rom_data[826]=16'b0111011101001111;
    rom_data[827]=16'b0011111011101010;
    rom_data[828]=16'b0111011101111000;
    rom_data[829]=16'b0011111111101000;
    rom_data[830]=16'b0111011110100001;
    rom_data[831]=16'b0100000011101010;
    rom_data[832]=16'b0111011111001001;
    rom_data[833]=16'b0100000111101110;
    rom_data[834]=16'b0111011111110010;
    rom_data[835]=16'b0100001011110110;
    rom_data[836]=16'b0111100000011010;
    rom_data[837]=16'b0100010000000001;
    rom_data[838]=16'b0111100001000010;
    rom_data[839]=16'b0100010100001111;
    rom_data[840]=16'b0111100001101010;
    rom_data[841]=16'b0100011000011111;
    rom_data[842]=16'b0111100010010001;
    rom_data[843]=16'b0100011100110001;
    rom_data[844]=16'b0111100010111000;
    rom_data[845]=16'b0100100001000110;
    rom_data[846]=16'b0111100011100000;
    rom_data[847]=16'b0100100101011100;
    rom_data[848]=16'b0111100100000111;
    rom_data[849]=16'b0100101001110101;
    rom_data[850]=16'b0111100100101101;
    rom_data[851]=16'b0100101110001111;
    rom_data[852]=16'b0111100101010100;
    rom_data[853]=16'b0100110010101011;
    rom_data[854]=16'b0111100101111011;
    rom_data[855]=16'b0100110111001001;
    rom_data[856]=16'b0111100110100001;
    rom_data[857]=16'b0100111011100111;
    rom_data[858]=16'b0111100111001000;
    rom_data[859]=16'b0101000000000111;
    rom_data[860]=16'b0111100111101110;
    rom_data[861]=16'b0101000100101000;
    rom_data[862]=16'b0111101000010100;
    rom_data[863]=16'b0101001001001011;
    rom_data[864]=16'b0111101000111010;
    rom_data[865]=16'b0101001101101110;
    rom_data[866]=16'b0111101001100000;
    rom_data[867]=16'b0101010010010001;
    rom_data[868]=16'b0111101010000110;
    rom_data[869]=16'b0101010110110110;
    rom_data[870]=16'b0111101010101100;
    rom_data[871]=16'b0101011011011011;
    rom_data[872]=16'b0111101011010010;
    rom_data[873]=16'b0101100000000000;
    rom_data[874]=16'b0111101011111000;
    rom_data[875]=16'b0101100100100110;
    rom_data[876]=16'b0111101100011110;
    rom_data[877]=16'b0101101001001101;
    rom_data[878]=16'b0111101101000100;
    rom_data[879]=16'b0101101101110011;
    rom_data[880]=16'b0111101101101010;
    rom_data[881]=16'b0101110010011010;
    rom_data[882]=16'b0111101110010000;
    rom_data[883]=16'b0101110111000001;
    rom_data[884]=16'b0111101110110111;
    rom_data[885]=16'b0101111011100111;
    rom_data[886]=16'b0111101111011101;
    rom_data[887]=16'b0110000000001110;
    rom_data[888]=16'b0111110000000011;
    rom_data[889]=16'b0110000100110100;
    rom_data[890]=16'b0111110000101001;
    rom_data[891]=16'b0110001001011010;
    rom_data[892]=16'b0111110001010000;
    rom_data[893]=16'b0110001110000000;
    rom_data[894]=16'b0111110001110110;
    rom_data[895]=16'b0110010010100101;
    rom_data[896]=16'b0111110010011101;
    rom_data[897]=16'b0110010111001001;
    rom_data[898]=16'b0111110011000100;
    rom_data[899]=16'b0110011011101101;
    rom_data[900]=16'b0111110011101011;
    rom_data[901]=16'b0110100000010000;
    rom_data[902]=16'b0111110100010010;
    rom_data[903]=16'b0110100100110010;
    rom_data[904]=16'b0111110100111001;
    rom_data[905]=16'b0110101001010011;
    rom_data[906]=16'b0111110101100001;
    rom_data[907]=16'b0110101101110100;
    rom_data[908]=16'b0111110110001001;
    rom_data[909]=16'b0110110010010010;
    rom_data[910]=16'b0111110110110001;
    rom_data[911]=16'b0110110110110000;
    rom_data[912]=16'b0111110111011001;
    rom_data[913]=16'b0110111011001100;
    rom_data[914]=16'b0111111000000001;
    rom_data[915]=16'b0110111111100111;
    rom_data[916]=16'b0111111000101010;
    rom_data[917]=16'b0111000100000000;
    rom_data[918]=16'b0111111001010011;
    rom_data[919]=16'b0111001000010111;
    rom_data[920]=16'b0111111001111100;
    rom_data[921]=16'b0111001100101100;
    rom_data[922]=16'b0111111010100101;
    rom_data[923]=16'b0111010000111111;
    rom_data[924]=16'b0111111011001111;
    rom_data[925]=16'b0111010101010000;
    rom_data[926]=16'b0111111011111001;
    rom_data[927]=16'b0111011001011111;
    rom_data[928]=16'b0111111100100100;
    rom_data[929]=16'b0111011101101010;
    rom_data[930]=16'b0111111101001111;
    rom_data[931]=16'b0111100001110011;
    rom_data[932]=16'b0111111101111010;
    rom_data[933]=16'b0111100101111010;
    rom_data[934]=16'b0111111110100110;
    rom_data[935]=16'b0111101001111101;
    rom_data[936]=16'b0111111111010010;
    rom_data[937]=16'b0111101101111100;
    rom_data[938]=16'b0111111111111110;
    rom_data[939]=16'b0111110001111000;
    rom_data[940]=16'b1000000000101011;
    rom_data[941]=16'b0111110101110000;
    rom_data[942]=16'b1000000001011001;
    rom_data[943]=16'b0111111001100100;
    rom_data[944]=16'b1000000010000110;
    rom_data[945]=16'b0111111101010100;
    rom_data[946]=16'b1000000010110101;
    rom_data[947]=16'b1000000000111111;
    rom_data[948]=16'b1000000011100100;
    rom_data[949]=16'b1000000100100101;
    rom_data[950]=16'b1000000100010011;
    rom_data[951]=16'b1000001000000101;
    rom_data[952]=16'b1000000101000011;
    rom_data[953]=16'b1000001011100000;
    rom_data[954]=16'b1000000101110011;
    rom_data[955]=16'b1000001110110101;
    rom_data[956]=16'b1000000110100100;
    rom_data[957]=16'b1000010010000100;
    rom_data[958]=16'b1000000111010101;
    rom_data[959]=16'b1000010101001100;
    rom_data[960]=16'b1000001000000111;
    rom_data[961]=16'b1000011000001100;
    rom_data[962]=16'b1000001000111010;
    rom_data[963]=16'b1000011011000101;
    rom_data[964]=16'b1000001001101101;
    rom_data[965]=16'b1000011101110101;
    rom_data[966]=16'b1000001010100000;
    rom_data[967]=16'b1000100000011101;
    rom_data[968]=16'b1000001011010100;
    rom_data[969]=16'b1000100010111011;
    rom_data[970]=16'b1000001100001000;
    rom_data[971]=16'b1000100101010000;
    rom_data[972]=16'b1000001100111101;
    rom_data[973]=16'b1000100111011010;
    rom_data[974]=16'b1000001101110001;
    rom_data[975]=16'b1000101001011010;
    rom_data[976]=16'b1000001110100111;
    rom_data[977]=16'b1000101011001110;
    rom_data[978]=16'b1000001111011100;
    rom_data[979]=16'b1000101100110110;
    rom_data[980]=16'b1000010000000010;
    rom_data[981]=16'b1000101110010010;
    rom_data[982]=16'b1000010000110111;
    rom_data[983]=16'b1000101111100010;
    rom_data[984]=16'b1000010001101100;
    rom_data[985]=16'b1000110000100100;
    rom_data[986]=16'b1000010010100001;
    rom_data[987]=16'b1000110001011000;
    rom_data[988]=16'b1000010011010101;
    rom_data[989]=16'b1000110001111110;
    rom_data[990]=16'b1000010100001010;
    rom_data[991]=16'b1000110010010110;
    rom_data[992]=16'b1000010100111110;
    rom_data[993]=16'b1000110010100000;
    rom_data[994]=16'b1000010101110010;
    rom_data[995]=16'b1000110010011011;
    rom_data[996]=16'b1000010110100110;
    rom_data[997]=16'b1000110010001000;
    rom_data[998]=16'b1000010111011001;
    rom_data[999]=16'b1000110001100110;
    rom_data[1000]=16'b1000011000001100;
    rom_data[1001]=16'b1000110000110110;
    rom_data[1002]=16'b1000011000111110;
    rom_data[1003]=16'b1000101111111001;
    rom_data[1004]=16'b1000011001110000;
    rom_data[1005]=16'b1000101110101101;
    rom_data[1006]=16'b1000011010100001;
    rom_data[1007]=16'b1000101101010101;
    rom_data[1008]=16'b1000011011010010;
    rom_data[1009]=16'b1000101011110000;
    rom_data[1010]=16'b1000011100000010;
    rom_data[1011]=16'b1000101001111110;
    rom_data[1012]=16'b1000011100110001;
    rom_data[1013]=16'b1000101000000000;
    rom_data[1014]=16'b1000011101100000;
    rom_data[1015]=16'b1000100101111000;
    rom_data[1016]=16'b1000011110001110;
    rom_data[1017]=16'b1000100011100100;
    rom_data[1018]=16'b1000011110111100;
    rom_data[1019]=16'b1000100001000111;
    rom_data[1020]=16'b1000011111101001;
    rom_data[1021]=16'b1000011110100000;
    rom_data[1022]=16'b1000100000010101;
    rom_data[1023]=16'b1000011011110000;
    rom_data[1024]=16'b1000100001000001;
    rom_data[1025]=16'b1000011000110111;
    rom_data[1026]=16'b1000100001101100;
    rom_data[1027]=16'b1000010101110110;
    rom_data[1028]=16'b1000100010010111;
    rom_data[1029]=16'b1000010010101110;
    rom_data[1030]=16'b1000100011000001;
    rom_data[1031]=16'b1000001111011110;
    rom_data[1032]=16'b1000100011101010;
    rom_data[1033]=16'b1000001100001000;
    rom_data[1034]=16'b1000100100010011;
    rom_data[1035]=16'b1000001000101100;
    rom_data[1036]=16'b1000100100111011;
    rom_data[1037]=16'b1000000101001010;
    rom_data[1038]=16'b1000100101100011;
    rom_data[1039]=16'b1000000001100011;
    rom_data[1040]=16'b1000100110001011;
    rom_data[1041]=16'b0111111101110110;
    rom_data[1042]=16'b1000100110110001;
    rom_data[1043]=16'b0111111010000101;
    rom_data[1044]=16'b1000100111011000;
    rom_data[1045]=16'b0111110110001111;
    rom_data[1046]=16'b1000100111111101;
    rom_data[1047]=16'b0111110010010101;
    rom_data[1048]=16'b1000101000100010;
    rom_data[1049]=16'b0111101110011000;
    rom_data[1050]=16'b1000101001000111;
    rom_data[1051]=16'b0111101010010110;
    rom_data[1052]=16'b1000101001101011;
    rom_data[1053]=16'b0111100110010010;
    rom_data[1054]=16'b1000101010001111;
    rom_data[1055]=16'b0111100010001010;
    rom_data[1056]=16'b1000101010110010;
    rom_data[1057]=16'b0111011101111111;
    rom_data[1058]=16'b1000101011010100;
    rom_data[1059]=16'b0111011001110001;
    rom_data[1060]=16'b1000101011110110;
    rom_data[1061]=16'b0111010101100001;
    rom_data[1062]=16'b1000101100011000;
    rom_data[1063]=16'b0111010001001111;
    rom_data[1064]=16'b1000101100111001;
    rom_data[1065]=16'b0111001100111010;
    rom_data[1066]=16'b1000101101011001;
    rom_data[1067]=16'b0111001000100011;
    rom_data[1068]=16'b1000101101111000;
    rom_data[1069]=16'b0111000100001011;
    rom_data[1070]=16'b1000101110010111;
    rom_data[1071]=16'b0110111111110001;
    rom_data[1072]=16'b1000101110110110;
    rom_data[1073]=16'b0110111011010101;
    rom_data[1074]=16'b1000101111010011;
    rom_data[1075]=16'b0110110110110111;
    rom_data[1076]=16'b1000101111110000;
    rom_data[1077]=16'b0110110010011000;
    rom_data[1078]=16'b1000110000001100;
    rom_data[1079]=16'b0110101101111000;
    rom_data[1080]=16'b1000110000100111;
    rom_data[1081]=16'b0110101001010111;
    rom_data[1082]=16'b1000110001000001;
    rom_data[1083]=16'b0110100100110101;
    rom_data[1084]=16'b1000110001011011;
    rom_data[1085]=16'b0110100000010010;
    rom_data[1086]=16'b1000110001110011;
    rom_data[1087]=16'b0110011011101111;
    rom_data[1088]=16'b1000110010001010;
    rom_data[1089]=16'b0110010111001010;
    rom_data[1090]=16'b1000110010100000;
    rom_data[1091]=16'b0110010010100101;
    rom_data[1092]=16'b1000110010100000;
    rom_data[1093]=16'b0110001101111111;
    rom_data[1094]=16'b1000110010001010;
    rom_data[1095]=16'b0110001001011001;
    rom_data[1096]=16'b1000110001110011;
    rom_data[1097]=16'b0110000100110011;
    rom_data[1098]=16'b1000110001011011;
    rom_data[1099]=16'b0110000000001101;
    rom_data[1100]=16'b1000110001000001;
    rom_data[1101]=16'b0101111011100110;
    rom_data[1102]=16'b1000110000100111;
    rom_data[1103]=16'b0101110110111111;
    rom_data[1104]=16'b1000110000001100;
    rom_data[1105]=16'b0101110010011001;
    rom_data[1106]=16'b1000101111110000;
    rom_data[1107]=16'b0101101101110010;
    rom_data[1108]=16'b1000101111010011;
    rom_data[1109]=16'b0101101001001100;
    rom_data[1110]=16'b1000101110110110;
    rom_data[1111]=16'b0101100100100110;
    rom_data[1112]=16'b1000101110010111;
    rom_data[1113]=16'b0101100000000000;
    rom_data[1114]=16'b1000101101111000;
    rom_data[1115]=16'b0101011011011011;
    rom_data[1116]=16'b1000101101011001;
    rom_data[1117]=16'b0101010110110111;
    rom_data[1118]=16'b1000101100111001;
    rom_data[1119]=16'b0101010010010011;
    rom_data[1120]=16'b1000101100011000;
    rom_data[1121]=16'b0101001101110000;
    rom_data[1122]=16'b1000101011110110;
    rom_data[1123]=16'b0101001001001110;
    rom_data[1124]=16'b1000101011010100;
    rom_data[1125]=16'b0101000100101100;
    rom_data[1126]=16'b1000101010110010;
    rom_data[1127]=16'b0101000000001100;
    rom_data[1128]=16'b1000101010001111;
    rom_data[1129]=16'b0100111011101101;
    rom_data[1130]=16'b1000101001101011;
    rom_data[1131]=16'b0100110111010000;
    rom_data[1132]=16'b1000101001000111;
    rom_data[1133]=16'b0100110010110100;
    rom_data[1134]=16'b1000101000100010;
    rom_data[1135]=16'b0100101110011001;
    rom_data[1136]=16'b1000100111111101;
    rom_data[1137]=16'b0100101010000000;
    rom_data[1138]=16'b1000100111011000;
    rom_data[1139]=16'b0100100101101001;
    rom_data[1140]=16'b1000100110110001;
    rom_data[1141]=16'b0100100001010100;
    rom_data[1142]=16'b1000100110001011;
    rom_data[1143]=16'b0100011101000001;
    rom_data[1144]=16'b1000100101100011;
    rom_data[1145]=16'b0100011000110000;
    rom_data[1146]=16'b1000100100111011;
    rom_data[1147]=16'b0100010100100001;
    rom_data[1148]=16'b1000100100010011;
    rom_data[1149]=16'b0100010000010101;
    rom_data[1150]=16'b1000100011101010;
    rom_data[1151]=16'b0100001100001100;
    rom_data[1152]=16'b1000100011000001;
    rom_data[1153]=16'b0100001000000110;
    rom_data[1154]=16'b1000100010010111;
    rom_data[1155]=16'b0100000100000011;
    rom_data[1156]=16'b1000100001101100;
    rom_data[1157]=16'b0100000000000100;
    rom_data[1158]=16'b1000100001000001;
    rom_data[1159]=16'b0011111100001000;
    rom_data[1160]=16'b1000100000010101;
    rom_data[1161]=16'b0011111000010000;
    rom_data[1162]=16'b1000011111101001;
    rom_data[1163]=16'b0011110100011100;
    rom_data[1164]=16'b1000011110111100;
    rom_data[1165]=16'b0011110000101100;
    rom_data[1166]=16'b1000011110001110;
    rom_data[1167]=16'b0011101101000001;
    rom_data[1168]=16'b1000011101100000;
    rom_data[1169]=16'b0011101001011011;
    rom_data[1170]=16'b1000011100110001;
    rom_data[1171]=16'b0011100101111010;
    rom_data[1172]=16'b1000011100000010;
    rom_data[1173]=16'b0011100010011111;
    rom_data[1174]=16'b1000011011010010;
    rom_data[1175]=16'b0011011111001010;
    rom_data[1176]=16'b1000011010100001;
    rom_data[1177]=16'b0011011011111100;
    rom_data[1178]=16'b1000011001110000;
    rom_data[1179]=16'b0011011000110100;
    rom_data[1180]=16'b1000011000111110;
    rom_data[1181]=16'b0011010101110100;
    rom_data[1182]=16'b1000011000001100;
    rom_data[1183]=16'b0011010010111011;
    rom_data[1184]=16'b1000010111011001;
    rom_data[1185]=16'b0011010000001011;
    rom_data[1186]=16'b1000010110100110;
    rom_data[1187]=16'b0011001101100011;
    rom_data[1188]=16'b1000010101110010;
    rom_data[1189]=16'b0011001011000101;
    rom_data[1190]=16'b1000010100111110;
    rom_data[1191]=16'b0011001000110000;
    rom_data[1192]=16'b1000010100001010;
    rom_data[1193]=16'b0011000110100110;
    rom_data[1194]=16'b1000010011010101;
    rom_data[1195]=16'b0011000100100110;
    rom_data[1196]=16'b1000010010100001;
    rom_data[1197]=16'b0011000010110010;
    rom_data[1198]=16'b1000010001101100;
    rom_data[1199]=16'b0011000001001001;
    rom_data[1200]=16'b1000010000110111;
    rom_data[1201]=16'b0010111111101101;
    rom_data[1202]=16'b1000010000000010;
    rom_data[1203]=16'b0010111110011110;
    rom_data[1204]=16'b1000001111011100;
    rom_data[1205]=16'b0010111101011100;
    rom_data[1206]=16'b1000001110100111;
    rom_data[1207]=16'b0010111100101000;
    rom_data[1208]=16'b1000001101110001;
    rom_data[1209]=16'b0010111100000010;
    rom_data[1210]=16'b1000001100111101;
    rom_data[1211]=16'b0010111011101010;
    rom_data[1212]=16'b1000001100001000;
    rom_data[1213]=16'b0010111011100000;
    rom_data[1214]=16'b1000001011010100;
    rom_data[1215]=16'b0010111011100101;
    rom_data[1216]=16'b1000001010100000;
    rom_data[1217]=16'b0010111011111000;
    rom_data[1218]=16'b1000001001101101;
    rom_data[1219]=16'b0010111100011010;
    rom_data[1220]=16'b1000001000111010;
    rom_data[1221]=16'b0010111101001010;
    rom_data[1222]=16'b1000001000000111;
    rom_data[1223]=16'b0010111110000111;
    rom_data[1224]=16'b1000000111010101;
    rom_data[1225]=16'b0010111111010011;
    rom_data[1226]=16'b1000000110100100;
    rom_data[1227]=16'b0011000000101011;
    rom_data[1228]=16'b1000000101110011;
    rom_data[1229]=16'b0011000010010001;
    rom_data[1230]=16'b1000000101000011;
    rom_data[1231]=16'b0011000100000010;
    rom_data[1232]=16'b1000000100010011;
    rom_data[1233]=16'b0011000110000000;
    rom_data[1234]=16'b1000000011100100;
    rom_data[1235]=16'b0011001000001000;
    rom_data[1236]=16'b1000000010110101;
    rom_data[1237]=16'b0011001010011100;
    rom_data[1238]=16'b1000000010000110;
    rom_data[1239]=16'b0011001100111001;
    rom_data[1240]=16'b1000000001011001;
    rom_data[1241]=16'b0011001111100000;
    rom_data[1242]=16'b1000000000101011;
    rom_data[1243]=16'b0011010010010001;
    rom_data[1244]=16'b0111111111111110;
    rom_data[1245]=16'b0011010101001001;
    rom_data[1246]=16'b0111111111010010;
    rom_data[1247]=16'b0011011000001010;
    rom_data[1248]=16'b0111111110100110;
    rom_data[1249]=16'b0011011011010010;
    rom_data[1250]=16'b0111111101111010;
    rom_data[1251]=16'b0011011110100010;
    rom_data[1252]=16'b0111111101001111;
    rom_data[1253]=16'b0011100001111000;
    rom_data[1254]=16'b0111111100100100;
    rom_data[1255]=16'b0011100101010100;
    rom_data[1256]=16'b0111111011111001;
    rom_data[1257]=16'b0011101000110110;
    rom_data[1258]=16'b0111111011001111;
    rom_data[1259]=16'b0011101100011101;
    rom_data[1260]=16'b0111111010100101;
    rom_data[1261]=16'b0011110000001010;
    rom_data[1262]=16'b0111111001111100;
    rom_data[1263]=16'b0011110011111011;
    rom_data[1264]=16'b0111111001010011;
    rom_data[1265]=16'b0011110111110001;
    rom_data[1266]=16'b0111111000101010;
    rom_data[1267]=16'b0011111011101011;
    rom_data[1268]=16'b0111111000000001;
    rom_data[1269]=16'b0011111111101001;
    rom_data[1270]=16'b0111110111011001;
    rom_data[1271]=16'b0100000011101010;
    rom_data[1272]=16'b0111110110110001;
    rom_data[1273]=16'b0100000111101111;
    rom_data[1274]=16'b0111110110001001;
    rom_data[1275]=16'b0100001011110110;
    rom_data[1276]=16'b0111110101100001;
    rom_data[1277]=16'b0100010000000001;
    rom_data[1278]=16'b0111110100111001;
    rom_data[1279]=16'b0100010100001111;
    rom_data[1280]=16'b0111110100010010;
    rom_data[1281]=16'b0100011000011111;
    rom_data[1282]=16'b0111110011101011;
    rom_data[1283]=16'b0100011100110001;
    rom_data[1284]=16'b0111110011000100;
    rom_data[1285]=16'b0100100001000110;
    rom_data[1286]=16'b0111110010011101;
    rom_data[1287]=16'b0100100101011101;
    rom_data[1288]=16'b0111110001110110;
    rom_data[1289]=16'b0100101001110101;
    rom_data[1290]=16'b0111110001010000;
    rom_data[1291]=16'b0100101110010000;
    rom_data[1292]=16'b0111110000101001;
    rom_data[1293]=16'b0100110010101100;
    rom_data[1294]=16'b0111110000000011;
    rom_data[1295]=16'b0100110111001001;
    rom_data[1296]=16'b0111101111011101;
    rom_data[1297]=16'b0100111011101000;
    rom_data[1298]=16'b0111101110110111;
    rom_data[1299]=16'b0101000000001000;
    rom_data[1300]=16'b0111101110010000;
    rom_data[1301]=16'b0101000100101001;
    rom_data[1302]=16'b0111101101101010;
    rom_data[1303]=16'b0101001001001011;
    rom_data[1304]=16'b0111101101000100;
    rom_data[1305]=16'b0101001101101110;
    rom_data[1306]=16'b0111101100011110;
    rom_data[1307]=16'b0101010010010010;
    rom_data[1308]=16'b0111101011111000;
    rom_data[1309]=16'b0101010110110110;
    rom_data[1310]=16'b0111101011010010;
    rom_data[1311]=16'b0101011011011011;
    rom_data[1312]=16'b0111101010101100;
    rom_data[1313]=16'b0101100000000001;
    rom_data[1314]=16'b0111101010000110;
    rom_data[1315]=16'b0101100100100111;
    rom_data[1316]=16'b0111101001100000;
    rom_data[1317]=16'b0101101001001101;
    rom_data[1318]=16'b0111101000111010;
    rom_data[1319]=16'b0101101101110100;
    rom_data[1320]=16'b0111101000010100;
    rom_data[1321]=16'b0101110010011010;
    rom_data[1322]=16'b0111100111101110;
    rom_data[1323]=16'b0101110111000001;
    rom_data[1324]=16'b0111100111001000;
    rom_data[1325]=16'b0101111011101000;
    rom_data[1326]=16'b0111100110100001;
    rom_data[1327]=16'b0110000000001110;
    rom_data[1328]=16'b0111100101111011;
    rom_data[1329]=16'b0110000100110100;
    rom_data[1330]=16'b0111100101010100;
    rom_data[1331]=16'b0110001001011010;
    rom_data[1332]=16'b0111100100101101;
    rom_data[1333]=16'b0110001110000000;
    rom_data[1334]=16'b0111100100000111;
    rom_data[1335]=16'b0110010010100101;
    rom_data[1336]=16'b0111100011100000;
    rom_data[1337]=16'b0110010111001010;
    rom_data[1338]=16'b0111100010111000;
    rom_data[1339]=16'b0110011011101101;
    rom_data[1340]=16'b0111100010010001;
    rom_data[1341]=16'b0110100000010000;
    rom_data[1342]=16'b0111100001101010;
    rom_data[1343]=16'b0110100100110011;
    rom_data[1344]=16'b0111100001000010;
    rom_data[1345]=16'b0110101001010100;
    rom_data[1346]=16'b0111100000011010;
    rom_data[1347]=16'b0110101101110100;
    rom_data[1348]=16'b0111011111110010;
    rom_data[1349]=16'b0110110010010011;
    rom_data[1350]=16'b0111011111001001;
    rom_data[1351]=16'b0110110110110000;
    rom_data[1352]=16'b0111011110100001;
    rom_data[1353]=16'b0110111011001101;
    rom_data[1354]=16'b0111011101111000;
    rom_data[1355]=16'b0110111111100111;
    rom_data[1356]=16'b0111011101001111;
    rom_data[1357]=16'b0111000100000000;
    rom_data[1358]=16'b0111011100100101;
    rom_data[1359]=16'b0111001000010111;
    rom_data[1360]=16'b0111011011111011;
    rom_data[1361]=16'b0111001100101100;
    rom_data[1362]=16'b0111011011010001;
    rom_data[1363]=16'b0111010001000000;
    rom_data[1364]=16'b0111011010100110;
    rom_data[1365]=16'b0111010101010000;
    rom_data[1366]=16'b0111011001111100;
    rom_data[1367]=16'b0111011001011111;
    rom_data[1368]=16'b0111011001010000;
    rom_data[1369]=16'b0111011101101011;
    rom_data[1370]=16'b0111011000100100;
    rom_data[1371]=16'b0111100001110100;
    rom_data[1372]=16'b0111010111111000;
    rom_data[1373]=16'b0111100101111010;
    rom_data[1374]=16'b0111010111001100;
    rom_data[1375]=16'b0111101001111101;
    rom_data[1376]=16'b0111010110011111;
    rom_data[1377]=16'b0111101101111100;
    rom_data[1378]=16'b0111010101110001;
    rom_data[1379]=16'b0111110001111000;
    rom_data[1380]=16'b0111010101000011;
    rom_data[1381]=16'b0111110101110001;
    rom_data[1382]=16'b0111010100010101;
    rom_data[1383]=16'b0111111001100101;
    rom_data[1384]=16'b0111010011100110;
    rom_data[1385]=16'b0111111101010100;
    rom_data[1386]=16'b0111010010110111;
    rom_data[1387]=16'b1000000000111111;
    rom_data[1388]=16'b0111010010000111;
    rom_data[1389]=16'b1000000100100101;
    rom_data[1390]=16'b0111010001010110;
    rom_data[1391]=16'b1000001000000110;
    rom_data[1392]=16'b0111010000100101;
    rom_data[1393]=16'b1000001011100001;
    rom_data[1394]=16'b0111001111110100;
    rom_data[1395]=16'b1000001110110110;
    rom_data[1396]=16'b0111001111000010;
    rom_data[1397]=16'b1000010010000100;
    rom_data[1398]=16'b0111001110001111;
    rom_data[1399]=16'b1000010101001100;
    rom_data[1400]=16'b0111001101011100;
    rom_data[1401]=16'b1000011000001100;
    rom_data[1402]=16'b0111001100101000;
    rom_data[1403]=16'b1000011011000101;
    rom_data[1404]=16'b0111001011110101;
    rom_data[1405]=16'b1000011101110101;
    rom_data[1406]=16'b0111001011000000;
    rom_data[1407]=16'b1000100000011101;
    rom_data[1408]=16'b0111001010001100;
    rom_data[1409]=16'b1000100010111011;
    rom_data[1410]=16'b0111001001010111;
    rom_data[1411]=16'b1000100101010000;
    rom_data[1412]=16'b0111001000100001;
    rom_data[1413]=16'b1000100111011010;
    rom_data[1414]=16'b0111000111101100;
    rom_data[1415]=16'b1000101001011010;
    rom_data[1416]=16'b0111000110110110;
    rom_data[1417]=16'b1000101011001110;
    rom_data[1418]=16'b0111000110000000;
    rom_data[1419]=16'b1000101100110111;
    rom_data[1420]=16'b0111000101001011;
    rom_data[1421]=16'b1000101110010011;
    rom_data[1422]=16'b0111000100010101;
    rom_data[1423]=16'b1000101111100010;
    rom_data[1424]=16'b0111000011011111;
    rom_data[1425]=16'b1000110000100100;
    rom_data[1426]=16'b0111000010101010;
    rom_data[1427]=16'b1000110001011000;
    rom_data[1428]=16'b0111000001110101;
    rom_data[1429]=16'b1000110001111110;
    rom_data[1430]=16'b0111000001000000;
    rom_data[1431]=16'b1000110010010110;
    rom_data[1432]=16'b0111000000001011;
    rom_data[1433]=16'b1000110010100000;
    rom_data[1434]=16'b0110111111010111;
    rom_data[1435]=16'b1000110010011011;
    rom_data[1436]=16'b0110111110100011;
    rom_data[1437]=16'b1000110010001000;
    rom_data[1438]=16'b0110111101110000;
    rom_data[1439]=16'b1000110001100110;
    rom_data[1440]=16'b0110111100111101;
    rom_data[1441]=16'b1000110000110110;
    rom_data[1442]=16'b0110111100001011;
    rom_data[1443]=16'b1000101111111001;
    rom_data[1444]=16'b0110111011011001;
    rom_data[1445]=16'b1000101110101101;
    rom_data[1446]=16'b0110111010100111;
    rom_data[1447]=16'b1000101101010101;
    rom_data[1448]=16'b0110111001110111;
    rom_data[1449]=16'b1000101011101111;
    rom_data[1450]=16'b0110111001000110;
    rom_data[1451]=16'b1000101001111110;
    rom_data[1452]=16'b0110111000010110;
    rom_data[1453]=16'b1000101000000000;
    rom_data[1454]=16'b0110110111100111;
    rom_data[1455]=16'b1000100101111000;
    rom_data[1456]=16'b0110110110111000;
    rom_data[1457]=16'b1000100011100100;
    rom_data[1458]=16'b0110110110001010;
    rom_data[1459]=16'b1000100001000111;
    rom_data[1460]=16'b0110110101011100;
    rom_data[1461]=16'b1000011110100000;
    rom_data[1462]=16'b0110110100101111;
    rom_data[1463]=16'b1000011011101111;
    rom_data[1464]=16'b0110110100000010;
    rom_data[1465]=16'b1000011000110111;
    rom_data[1466]=16'b0110110011010101;
    rom_data[1467]=16'b1000010101110110;
    rom_data[1468]=16'b0110110010101001;
    rom_data[1469]=16'b1000010010101110;
    rom_data[1470]=16'b0110110001111101;
    rom_data[1471]=16'b1000001111011110;
    rom_data[1472]=16'b0110110001010010;
    rom_data[1473]=16'b1000001100001000;
    rom_data[1474]=16'b0110110000100111;
    rom_data[1475]=16'b1000001000101100;
    rom_data[1476]=16'b0110101111111101;
    rom_data[1477]=16'b1000000101001010;
    rom_data[1478]=16'b0110101111010011;
    rom_data[1479]=16'b1000000001100010;
    rom_data[1480]=16'b0110101110101001;
    rom_data[1481]=16'b0111111101110110;
    rom_data[1482]=16'b0110101101111111;
    rom_data[1483]=16'b0111111010000101;
    rom_data[1484]=16'b0110101101010110;
    rom_data[1485]=16'b0111110110001111;
    rom_data[1486]=16'b0110101100101101;
    rom_data[1487]=16'b0111110010010101;
    rom_data[1488]=16'b0110101100000100;
    rom_data[1489]=16'b0111101110010111;
    rom_data[1490]=16'b0110101011011100;
    rom_data[1491]=16'b0111101010010110;
    rom_data[1492]=16'b0110101010110100;
    rom_data[1493]=16'b0111100110010001;
    rom_data[1494]=16'b0110101010001100;
    rom_data[1495]=16'b0111100010001001;
    rom_data[1496]=16'b0110101001100100;
    rom_data[1497]=16'b0111011101111111;
    rom_data[1498]=16'b0110101000111101;
    rom_data[1499]=16'b0111011001110001;
    rom_data[1500]=16'b0110101000010110;
    rom_data[1501]=16'b0111010101100001;
    rom_data[1502]=16'b0110100111101110;
    rom_data[1503]=16'b0111010001001110;
    rom_data[1504]=16'b0110100111000111;
    rom_data[1505]=16'b0111001100111010;
    rom_data[1506]=16'b0110100110100001;
    rom_data[1507]=16'b0111001000100011;
    rom_data[1508]=16'b0110100101111010;
    rom_data[1509]=16'b0111000100001011;
    rom_data[1510]=16'b0110100101010011;
    rom_data[1511]=16'b0110111111110000;
    rom_data[1512]=16'b0110100100101101;
    rom_data[1513]=16'b0110111011010100;
    rom_data[1514]=16'b0110100100000110;
    rom_data[1515]=16'b0110110110110111;
    rom_data[1516]=16'b0110100011100000;
    rom_data[1517]=16'b0110110010011000;
    rom_data[1518]=16'b0110100010111010;
    rom_data[1519]=16'b0110101101111000;
    rom_data[1520]=16'b0110100010010100;
    rom_data[1521]=16'b0110101001010111;
    rom_data[1522]=16'b0110100001101110;
    rom_data[1523]=16'b0110100100110101;
    rom_data[1524]=16'b0110100001001000;
    rom_data[1525]=16'b0110100000010010;
    rom_data[1526]=16'b0110100000100010;
    rom_data[1527]=16'b0110011011101110;
    rom_data[1528]=16'b0110011111111100;
    rom_data[1529]=16'b0110010111001010;
    rom_data[1530]=16'b0110011111010110;
    rom_data[1531]=16'b0110010010100101;
    rom_data[1532]=16'b0110011110110000;
    rom_data[1533]=16'b0110001101111111;
    rom_data[1534]=16'b0110011110001010;
    rom_data[1535]=16'b0110001001011001;
    rom_data[1536]=16'b0110011101100100;
    rom_data[1537]=16'b0110000100110011;
    rom_data[1538]=16'b0110011100111110;
    rom_data[1539]=16'b0110000000001100;
    rom_data[1540]=16'b0110011100010111;
    rom_data[1541]=16'b0101111011100110;
    rom_data[1542]=16'b0110011011110001;
    rom_data[1543]=16'b0101110110111111;
    rom_data[1544]=16'b0110011011001011;
    rom_data[1545]=16'b0101110010011000;
    rom_data[1546]=16'b0110011010100101;
    rom_data[1547]=16'b0101101101110010;
    rom_data[1548]=16'b0110011001111110;
    rom_data[1549]=16'b0101101001001011;
    rom_data[1550]=16'b0110011001011000;
    rom_data[1551]=16'b0101100100100101;
    rom_data[1552]=16'b0110011000110001;
    rom_data[1553]=16'b0101100000000000;
    rom_data[1554]=16'b0110011000001010;
    rom_data[1555]=16'b0101011011011011;
    rom_data[1556]=16'b0110010111100011;
    rom_data[1557]=16'b0101010110110110;
    rom_data[1558]=16'b0110010110111100;
    rom_data[1559]=16'b0101010010010010;
    rom_data[1560]=16'b0110010110010101;
    rom_data[1561]=16'b0101001101101111;
    rom_data[1562]=16'b0110010101101101;
    rom_data[1563]=16'b0101001001001101;
    rom_data[1564]=16'b0110010101000101;
    rom_data[1565]=16'b0101000100101100;
    rom_data[1566]=16'b0110010100011101;
    rom_data[1567]=16'b0101000000001100;
    rom_data[1568]=16'b0110010011110101;
    rom_data[1569]=16'b0100111011101101;
    rom_data[1570]=16'b0110010011001101;
    rom_data[1571]=16'b0100110111001111;
    rom_data[1572]=16'b0110010010100100;
    rom_data[1573]=16'b0100110010110011;
    rom_data[1574]=16'b0110010001111011;
    rom_data[1575]=16'b0100101110011001;
    rom_data[1576]=16'b0110010001010010;
    rom_data[1577]=16'b0100101010000000;
    rom_data[1578]=16'b0110010000101000;
    rom_data[1579]=16'b0100100101101001;
    rom_data[1580]=16'b0110001111111111;
    rom_data[1581]=16'b0100100001010011;
    rom_data[1582]=16'b0110001111010100;
    rom_data[1583]=16'b0100011101000000;
    rom_data[1584]=16'b0110001110101010;
    rom_data[1585]=16'b0100011000101111;
    rom_data[1586]=16'b0110001101111111;
    rom_data[1587]=16'b0100010100100001;
    rom_data[1588]=16'b0110001101010100;
    rom_data[1589]=16'b0100010000010101;
    rom_data[1590]=16'b0110001100101000;
    rom_data[1591]=16'b0100001100001100;
    rom_data[1592]=16'b0110001011111100;
    rom_data[1593]=16'b0100001000000110;
    rom_data[1594]=16'b0110001011001111;
    rom_data[1595]=16'b0100000100000011;
    rom_data[1596]=16'b0110001010100010;
    rom_data[1597]=16'b0100000000000011;
    rom_data[1598]=16'b0110001001110101;
    rom_data[1599]=16'b0011111100000111;
    rom_data[1600]=16'b0110001001000111;
    rom_data[1601]=16'b0011111000001111;
    rom_data[1602]=16'b0110001000011000;
    rom_data[1603]=16'b0011110100011011;
    rom_data[1604]=16'b0110000111101001;
    rom_data[1605]=16'b0011110000101100;
    rom_data[1606]=16'b0110000110111010;
    rom_data[1607]=16'b0011101101000001;
    rom_data[1608]=16'b0110000110001010;
    rom_data[1609]=16'b0011101001011011;
    rom_data[1610]=16'b0110000101011010;
    rom_data[1611]=16'b0011100101111010;
    rom_data[1612]=16'b0110000100101001;
    rom_data[1613]=16'b0011100010011111;
    rom_data[1614]=16'b0110000011110111;
    rom_data[1615]=16'b0011011111001010;
    rom_data[1616]=16'b0110000011000101;
    rom_data[1617]=16'b0011011011111100;
    rom_data[1618]=16'b0110000010010010;
    rom_data[1619]=16'b0011011000110100;
    rom_data[1620]=16'b0110000001011111;
    rom_data[1621]=16'b0011010101110100;
    rom_data[1622]=16'b0110000000101100;
    rom_data[1623]=16'b0011010010111011;
    rom_data[1624]=16'b0101111111111000;
    rom_data[1625]=16'b0011010000001011;
    rom_data[1626]=16'b0101111111000100;
    rom_data[1627]=16'b0011001101100011;
    rom_data[1628]=16'b0101111110001111;
    rom_data[1629]=16'b0011001011000101;
    rom_data[1630]=16'b0101111101011010;
    rom_data[1631]=16'b0011001000110000;
    rom_data[1632]=16'b0101111100100101;
    rom_data[1633]=16'b0011000110100110;
    rom_data[1634]=16'b0101111011101111;
    rom_data[1635]=16'b0011000100100110;
    rom_data[1636]=16'b0101111010111010;
    rom_data[1637]=16'b0011000010110010;
    rom_data[1638]=16'b0101111010000100;
    rom_data[1639]=16'b0011000001001001;
    rom_data[1640]=16'b0101111001001110;
    rom_data[1641]=16'b0010111111101101;
    rom_data[1642]=16'b0101111000011000;
    rom_data[1643]=16'b0010111110011110;
    rom_data[1644]=16'b0101110111100011;
    rom_data[1645]=16'b0010111101011100;
    rom_data[1646]=16'b0101110110101101;
    rom_data[1647]=16'b0010111100101000;
    rom_data[1648]=16'b0101110101111000;
    rom_data[1649]=16'b0010111100000010;
    rom_data[1650]=16'b0101110101000011;
    rom_data[1651]=16'b0010111011101010;
    rom_data[1652]=16'b0101110100001111;
    rom_data[1653]=16'b0010111011100000;
    rom_data[1654]=16'b0101110011011011;
    rom_data[1655]=16'b0010111011100101;
    rom_data[1656]=16'b0101110010100111;
    rom_data[1657]=16'b0010111011111000;
    rom_data[1658]=16'b0101110001110011;
    rom_data[1659]=16'b0010111100011010;
    rom_data[1660]=16'b0101110001000001;
    rom_data[1661]=16'b0010111101001010;
    rom_data[1662]=16'b0101110000001110;
    rom_data[1663]=16'b0010111110000111;
    rom_data[1664]=16'b0101101111011100;
    rom_data[1665]=16'b0010111111010011;
    rom_data[1666]=16'b0101101110101011;
    rom_data[1667]=16'b0011000000101011;
    rom_data[1668]=16'b0101101101111010;
    rom_data[1669]=16'b0011000010010001;
    rom_data[1670]=16'b0101101101001010;
    rom_data[1671]=16'b0011000100000010;
    rom_data[1672]=16'b0101101100011010;
    rom_data[1673]=16'b0011000110000000;
    rom_data[1674]=16'b0101101011101010;
    rom_data[1675]=16'b0011001000001000;
    rom_data[1676]=16'b0101101010111100;
    rom_data[1677]=16'b0011001010011100;
    rom_data[1678]=16'b0101101010001101;
    rom_data[1679]=16'b0011001100111001;
    rom_data[1680]=16'b0101101001011111;
    rom_data[1681]=16'b0011001111100001;
    rom_data[1682]=16'b0101101000110010;
    rom_data[1683]=16'b0011010010010001;
    rom_data[1684]=16'b0101101000000101;
    rom_data[1685]=16'b0011010101001010;
    rom_data[1686]=16'b0101100111011001;
    rom_data[1687]=16'b0011011000001010;
    rom_data[1688]=16'b0101100110101100;
    rom_data[1689]=16'b0011011011010011;
    rom_data[1690]=16'b0101100110000001;
    rom_data[1691]=16'b0011011110100010;
    rom_data[1692]=16'b0101100101010110;
    rom_data[1693]=16'b0011100001111000;
    rom_data[1694]=16'b0101100100101011;
    rom_data[1695]=16'b0011100101010100;
    rom_data[1696]=16'b0101100100000000;
    rom_data[1697]=16'b0011101000110110;
    rom_data[1698]=16'b0101100011010110;
    rom_data[1699]=16'b0011101100011110;
    rom_data[1700]=16'b0101100010101100;
    rom_data[1701]=16'b0011110000001010;
    rom_data[1702]=16'b0101100010000011;
    rom_data[1703]=16'b0011110011111011;
    rom_data[1704]=16'b0101100001011001;
    rom_data[1705]=16'b0011110111110001;
    rom_data[1706]=16'b0101100000110001;
    rom_data[1707]=16'b0011111011101011;
    rom_data[1708]=16'b0101100000001000;
    rom_data[1709]=16'b0011111111101001;
    rom_data[1710]=16'b0101011111100000;
    rom_data[1711]=16'b0100000011101010;
    rom_data[1712]=16'b0101011110110111;
    rom_data[1713]=16'b0100000111101111;
    rom_data[1714]=16'b0101011110001111;
    rom_data[1715]=16'b0100001011110111;
    rom_data[1716]=16'b0101011101101000;
    rom_data[1717]=16'b0100010000000010;
    rom_data[1718]=16'b0101011101000000;
    rom_data[1719]=16'b0100010100001111;
    rom_data[1720]=16'b0101011100011001;
    rom_data[1721]=16'b0100011000011111;
    rom_data[1722]=16'b0101011011110010;
    rom_data[1723]=16'b0100011100110010;
    rom_data[1724]=16'b0101011011001011;
    rom_data[1725]=16'b0100100001000110;
    rom_data[1726]=16'b0101011010100100;
    rom_data[1727]=16'b0100100101011101;
    rom_data[1728]=16'b0101011001111101;
    rom_data[1729]=16'b0100101001110110;
    rom_data[1730]=16'b0101011001010111;
    rom_data[1731]=16'b0100101110010000;
    rom_data[1732]=16'b0101011000110000;
    rom_data[1733]=16'b0100110010101100;
    rom_data[1734]=16'b0101011000001010;
    rom_data[1735]=16'b0100110111001001;
    rom_data[1736]=16'b0101010111100100;
    rom_data[1737]=16'b0100111011101000;
    rom_data[1738]=16'b0101010110111101;
    rom_data[1739]=16'b0101000000001000;
    rom_data[1740]=16'b0101010110010111;
    rom_data[1741]=16'b0101000100101001;
    rom_data[1742]=16'b0101010101110001;
    rom_data[1743]=16'b0101001001001011;
    rom_data[1744]=16'b0101010101001011;
    rom_data[1745]=16'b0101001101101110;
    rom_data[1746]=16'b0101010100100101;
    rom_data[1747]=16'b0101010010010010;
    rom_data[1748]=16'b0101010011111111;
    rom_data[1749]=16'b0101010110110110;
    rom_data[1750]=16'b0101010011011001;
    rom_data[1751]=16'b0101011011011100;
    rom_data[1752]=16'b0101010010110011;
    rom_data[1753]=16'b0101100000000001;
    rom_data[1754]=16'b0101010010001101;
    rom_data[1755]=16'b0101100100100111;
    rom_data[1756]=16'b0101010001100111;
    rom_data[1757]=16'b0101101001001101;
    rom_data[1758]=16'b0101010001000001;
    rom_data[1759]=16'b0101101101110100;
    rom_data[1760]=16'b0101010000011011;
    rom_data[1761]=16'b0101110010011011;
    rom_data[1762]=16'b0101001111110101;
    rom_data[1763]=16'b0101110111000001;
    rom_data[1764]=16'b0101001111001110;
    rom_data[1765]=16'b0101111011101000;
    rom_data[1766]=16'b0101001110101000;
    rom_data[1767]=16'b0110000000001110;
    rom_data[1768]=16'b0101001110000010;
    rom_data[1769]=16'b0110000100110101;
    rom_data[1770]=16'b0101001101011011;
    rom_data[1771]=16'b0110001001011011;
    rom_data[1772]=16'b0101001100110100;
    rom_data[1773]=16'b0110001110000000;
    rom_data[1774]=16'b0101001100001101;
    rom_data[1775]=16'b0110010010100101;
    rom_data[1776]=16'b0101001011100110;
    rom_data[1777]=16'b0110010111001010;
    rom_data[1778]=16'b0101001010111111;
    rom_data[1779]=16'b0110011011101110;
    rom_data[1780]=16'b0101001010011000;
    rom_data[1781]=16'b0110100000010001;
    rom_data[1782]=16'b0101001001110000;
    rom_data[1783]=16'b0110100100110011;
    rom_data[1784]=16'b0101001001001001;
    rom_data[1785]=16'b0110101001010100;
    rom_data[1786]=16'b0101001000100001;
    rom_data[1787]=16'b0110101101110100;
    rom_data[1788]=16'b0101000111111001;
    rom_data[1789]=16'b0110110010010011;
    rom_data[1790]=16'b0101000111010000;
    rom_data[1791]=16'b0110110110110001;
    rom_data[1792]=16'b0101000110101000;
    rom_data[1793]=16'b0110111011001101;
    rom_data[1794]=16'b0101000101111111;
    rom_data[1795]=16'b0110111111100111;
    rom_data[1796]=16'b0101000101010101;
    rom_data[1797]=16'b0111000100000000;
    rom_data[1798]=16'b0101000100101100;
    rom_data[1799]=16'b0111001000011000;
    rom_data[1800]=16'b0101000100000010;
    rom_data[1801]=16'b0111001100101101;
    rom_data[1802]=16'b0101000011011000;
    rom_data[1803]=16'b0111010001000000;
    rom_data[1804]=16'b0101000010101101;
    rom_data[1805]=16'b0111010101010001;
    rom_data[1806]=16'b0101000010000010;
    rom_data[1807]=16'b0111011001011111;
    rom_data[1808]=16'b0101000001010111;
    rom_data[1809]=16'b0111011101101011;
    rom_data[1810]=16'b0101000000101011;
    rom_data[1811]=16'b0111100001110100;
    rom_data[1812]=16'b0100111111111111;
    rom_data[1813]=16'b0111100101111010;
    rom_data[1814]=16'b0100111111010011;
    rom_data[1815]=16'b0111101001111101;
    rom_data[1816]=16'b0100111110100110;
    rom_data[1817]=16'b0111101101111101;
    rom_data[1818]=16'b0100111101111000;
    rom_data[1819]=16'b0111110001111001;
    rom_data[1820]=16'b0100111101001010;
    rom_data[1821]=16'b0111110101110001;
    rom_data[1822]=16'b0100111100011100;
    rom_data[1823]=16'b0111111001100101;
    rom_data[1824]=16'b0100111011101101;
    rom_data[1825]=16'b0111111101010100;
    rom_data[1826]=16'b0100111010111101;
    rom_data[1827]=16'b1000000000111111;
    rom_data[1828]=16'b0100111010001101;
    rom_data[1829]=16'b1000000100100101;
    rom_data[1830]=16'b0100111001011101;
    rom_data[1831]=16'b1000001000000110;
    rom_data[1832]=16'b0100111000101100;
    rom_data[1833]=16'b1000001011100001;
    rom_data[1834]=16'b0100110111111010;
    rom_data[1835]=16'b1000001110110110;
    rom_data[1836]=16'b0100110111001000;
    rom_data[1837]=16'b1000010010000100;
    rom_data[1838]=16'b0100110110010110;
    rom_data[1839]=16'b1000010101001100;
    rom_data[1840]=16'b0100110101100011;
    rom_data[1841]=16'b1000011000001100;
    rom_data[1842]=16'b0100110100101111;
    rom_data[1843]=16'b1000011011000101;
    rom_data[1844]=16'b0100110011111011;
    rom_data[1845]=16'b1000011101110101;
    rom_data[1846]=16'b0100110011000111;
    rom_data[1847]=16'b1000100000011101;
    rom_data[1848]=16'b0100110010010010;
    rom_data[1849]=16'b1000100010111011;
    rom_data[1850]=16'b0100110001011101;
    rom_data[1851]=16'b1000100101010000;
    rom_data[1852]=16'b0100110000101000;
    rom_data[1853]=16'b1000100111011011;
    rom_data[1854]=16'b0100101111110011;
    rom_data[1855]=16'b1000101001011010;
    rom_data[1856]=16'b0100101110111101;
    rom_data[1857]=16'b1000101011001110;
    rom_data[1858]=16'b0100101110000111;
    rom_data[1859]=16'b1000101100110111;
    rom_data[1860]=16'b0100101101010010;
    rom_data[1861]=16'b1000101110010011;
    rom_data[1862]=16'b0100101100011100;
    rom_data[1863]=16'b1000101111100010;
    rom_data[1864]=16'b0100101011100110;
    rom_data[1865]=16'b1000110000100100;
    rom_data[1866]=16'b0100101010110001;
    rom_data[1867]=16'b1000110001011000;
    rom_data[1868]=16'b0100101001111100;
    rom_data[1869]=16'b1000110001111110;
    rom_data[1870]=16'b0100101001000111;
    rom_data[1871]=16'b1000110010010110;
    rom_data[1872]=16'b0100101000010010;
    rom_data[1873]=16'b1000110010100000;
    rom_data[1874]=16'b0100100111011110;
    rom_data[1875]=16'b1000110010011011;
    rom_data[1876]=16'b0100100110101010;
    rom_data[1877]=16'b1000110010001000;
    rom_data[1878]=16'b0100100101110111;
    rom_data[1879]=16'b1000110001100110;
    rom_data[1880]=16'b0100100101000100;
    rom_data[1881]=16'b1000110000110110;
    rom_data[1882]=16'b0100100100010010;
    rom_data[1883]=16'b1000101111111001;
    rom_data[1884]=16'b0100100011100000;
    rom_data[1885]=16'b1000101110101101;
    rom_data[1886]=16'b0100100010101110;
    rom_data[1887]=16'b1000101101010101;
    rom_data[1888]=16'b0100100001111101;
    rom_data[1889]=16'b1000101011101111;
    rom_data[1890]=16'b0100100001001101;
    rom_data[1891]=16'b1000101001111110;
    rom_data[1892]=16'b0100100000011101;
    rom_data[1893]=16'b1000101000000000;
    rom_data[1894]=16'b0100011111101110;
    rom_data[1895]=16'b1000100101110111;
    rom_data[1896]=16'b0100011110111111;
    rom_data[1897]=16'b1000100011100100;
    rom_data[1898]=16'b0100011110010001;
    rom_data[1899]=16'b1000100001000110;
    rom_data[1900]=16'b0100011101100011;
    rom_data[1901]=16'b1000011110011111;
    rom_data[1902]=16'b0100011100110101;
    rom_data[1903]=16'b1000011011101111;
    rom_data[1904]=16'b0100011100001000;
    rom_data[1905]=16'b1000011000110110;
    rom_data[1906]=16'b0100011011011100;
    rom_data[1907]=16'b1000010101110110;
    rom_data[1908]=16'b0100011010110000;
    rom_data[1909]=16'b1000010010101101;
    rom_data[1910]=16'b0100011010000100;
    rom_data[1911]=16'b1000001111011110;
    rom_data[1912]=16'b0100011001011001;
    rom_data[1913]=16'b1000001100001000;
    rom_data[1914]=16'b0100011000101110;
    rom_data[1915]=16'b1000001000101100;
    rom_data[1916]=16'b0100011000000100;
    rom_data[1917]=16'b1000000101001010;
    rom_data[1918]=16'b0100010111011001;
    rom_data[1919]=16'b1000000001100010;
    rom_data[1920]=16'b0100010110110000;
    rom_data[1921]=16'b0111111101110110;
    rom_data[1922]=16'b0100010110000110;
    rom_data[1923]=16'b0111111010000100;
    rom_data[1924]=16'b0100010101011101;
    rom_data[1925]=16'b0111110110001111;
    rom_data[1926]=16'b0100010100110100;
    rom_data[1927]=16'b0111110010010101;
    rom_data[1928]=16'b0100010100001011;
    rom_data[1929]=16'b0111101110010111;
    rom_data[1930]=16'b0100010011100011;
    rom_data[1931]=16'b0111101010010110;
    rom_data[1932]=16'b0100010010111011;
    rom_data[1933]=16'b0111100110010001;
    rom_data[1934]=16'b0100010010010011;
    rom_data[1935]=16'b0111100010001001;
    rom_data[1936]=16'b0100010001101011;
    rom_data[1937]=16'b0111011101111110;
    rom_data[1938]=16'b0100010001000100;
    rom_data[1939]=16'b0111011001110001;
    rom_data[1940]=16'b0100010000011100;
    rom_data[1941]=16'b0111010101100001;
    rom_data[1942]=16'b0100001111110101;
    rom_data[1943]=16'b0111010001001110;
    rom_data[1944]=16'b0100001111001110;
    rom_data[1945]=16'b0111001100111010;
    rom_data[1946]=16'b0100001110100111;
    rom_data[1947]=16'b0111001000100011;
    rom_data[1948]=16'b0100001110000001;
    rom_data[1949]=16'b0111000100001010;
    rom_data[1950]=16'b0100001101011010;
    rom_data[1951]=16'b0110111111110000;
    rom_data[1952]=16'b0100001100110100;
    rom_data[1953]=16'b0110111011010100;
    rom_data[1954]=16'b0100001100001101;
    rom_data[1955]=16'b0110110110110111;
    rom_data[1956]=16'b0100001011100111;
    rom_data[1957]=16'b0110110010011000;
    rom_data[1958]=16'b0100001011000001;
    rom_data[1959]=16'b0110101101111000;
    rom_data[1960]=16'b0100001010011011;
    rom_data[1961]=16'b0110101001010111;
    rom_data[1962]=16'b0100001001110101;
    rom_data[1963]=16'b0110100100110101;
    rom_data[1964]=16'b0100001001001111;
    rom_data[1965]=16'b0110100000010010;
    rom_data[1966]=16'b0100001000101001;
    rom_data[1967]=16'b0110011011101110;
    rom_data[1968]=16'b0100001000000011;
    rom_data[1969]=16'b0110010111001001;
    rom_data[1970]=16'b0100000111011101;
    rom_data[1971]=16'b0110010010100100;
    rom_data[1972]=16'b0100000110110111;
    rom_data[1973]=16'b0110001101111111;
    rom_data[1974]=16'b0100000110010001;
    rom_data[1975]=16'b0110001001011001;
    rom_data[1976]=16'b0100000101101011;
    rom_data[1977]=16'b0110000100110010;
    rom_data[1978]=16'b0100000101000100;
    rom_data[1979]=16'b0110000000001100;
    rom_data[1980]=16'b0100000100011110;
    rom_data[1981]=16'b0101111011100101;
    rom_data[1982]=16'b0100000011111000;
    rom_data[1983]=16'b0101110110111111;
    rom_data[1984]=16'b0100000011010010;
    rom_data[1985]=16'b0101110010011000;
    rom_data[1986]=16'b0100000010101011;
    rom_data[1987]=16'b0101101101110001;
    rom_data[1988]=16'b0100000010000101;
    rom_data[1989]=16'b0101101001001011;
    rom_data[1990]=16'b0100000001011110;
    rom_data[1991]=16'b0101100100100101;
    rom_data[1992]=16'b0100000000111000;
    rom_data[1993]=16'b0101100000000000;
    rom_data[1994]=16'b0100000000010001;
    rom_data[1995]=16'b0101011011011010;
    rom_data[1996]=16'b0011111111101010;
    rom_data[1997]=16'b0101010110110110;
    rom_data[1998]=16'b0011111111000011;
    rom_data[1999]=16'b0101010010010010;
    rom_data[2000]=16'b0011111110011011;
    rom_data[2001]=16'b0101001101101111;
    rom_data[2002]=16'b0011111101110100;
    rom_data[2003]=16'b0101001001001101;
    rom_data[2004]=16'b0011111101001100;
    rom_data[2005]=16'b0101000100101100;
    rom_data[2006]=16'b0011111100100100;
    rom_data[2007]=16'b0101000000001100;
    rom_data[2008]=16'b0011111011111100;
    rom_data[2009]=16'b0100111011101101;
    rom_data[2010]=16'b0011111011010100;
    rom_data[2011]=16'b0100110111001111;
    rom_data[2012]=16'b0011111010101011;
    rom_data[2013]=16'b0100110010110011;
    rom_data[2014]=16'b0011111010000010;
    rom_data[2015]=16'b0100101110011000;
    rom_data[2016]=16'b0011111001011001;
    rom_data[2017]=16'b0100101001111111;
    rom_data[2018]=16'b0011111000101111;
    rom_data[2019]=16'b0100100101101000;
    rom_data[2020]=16'b0011111000000101;
    rom_data[2021]=16'b0100100001010011;
    rom_data[2022]=16'b0011110111011011;
    rom_data[2023]=16'b0100011101000000;
    rom_data[2024]=16'b0011110110110001;
    rom_data[2025]=16'b0100011000101111;
    rom_data[2026]=16'b0011110110000110;
    rom_data[2027]=16'b0100010100100001;
    rom_data[2028]=16'b0011110101011010;
    rom_data[2029]=16'b0100010000010101;
    rom_data[2030]=16'b0011110100101111;
    rom_data[2031]=16'b0100001100001100;
    rom_data[2032]=16'b0011110100000011;
    rom_data[2033]=16'b0100001000000110;
    rom_data[2034]=16'b0011110011010110;
    rom_data[2035]=16'b0100000100000011;
    rom_data[2036]=16'b0011110010101001;
    rom_data[2037]=16'b0100000000000011;
    rom_data[2038]=16'b0011110001111100;
    rom_data[2039]=16'b0011111100000111;
    rom_data[2040]=16'b0011110001001110;
    rom_data[2041]=16'b0011111000001111;
    rom_data[2042]=16'b0011110000011111;
    rom_data[2043]=16'b0011110100011011;
    rom_data[2044]=16'b0011101111110000;
    rom_data[2045]=16'b0011110000101011;
    rom_data[2046]=16'b0011101111000001;
    rom_data[2047]=16'b0011101101000001;
    rom_data[2048]=16'b0011101110010001;
    rom_data[2049]=16'b0011101001011011;
    rom_data[2050]=16'b0011101101100000;
    rom_data[2051]=16'b0011100101111010;
    rom_data[2052]=16'b0011101100101111;
    rom_data[2053]=16'b0011100010011111;
    rom_data[2054]=16'b0011101011111110;
    rom_data[2055]=16'b0011011111001010;
    rom_data[2056]=16'b0011101011001100;
    rom_data[2057]=16'b0011011011111100;
    rom_data[2058]=16'b0011101010011001;
    rom_data[2059]=16'b0011011000110100;
    rom_data[2060]=16'b0011101001100110;
    rom_data[2061]=16'b0011010101110100;
    rom_data[2062]=16'b0011101000110011;
    rom_data[2063]=16'b0011010010111011;
    rom_data[2064]=16'b0011100111111111;
    rom_data[2065]=16'b0011010000001011;
    rom_data[2066]=16'b0011100111001010;
    rom_data[2067]=16'b0011001101100011;
    rom_data[2068]=16'b0011100110010110;
    rom_data[2069]=16'b0011001011000100;
    rom_data[2070]=16'b0011100101100001;
    rom_data[2071]=16'b0011001000110000;
    rom_data[2072]=16'b0011100100101100;
    rom_data[2073]=16'b0011000110100101;
    rom_data[2074]=16'b0011100011110110;
    rom_data[2075]=16'b0011000100100110;
    rom_data[2076]=16'b0011100011000000;
    rom_data[2077]=16'b0011000010110010;
    rom_data[2078]=16'b0011100010001011;
    rom_data[2079]=16'b0011000001001001;
    rom_data[2080]=16'b0011100001010101;
    rom_data[2081]=16'b0010111111101101;
    rom_data[2082]=16'b0011100000110001;
    rom_data[2083]=16'b0010111110011110;
    rom_data[2084]=16'b0011011111111100;
    rom_data[2085]=16'b0010111101011100;
    rom_data[2086]=16'b0011011111001000;
    rom_data[2087]=16'b0010111100101000;
    rom_data[2088]=16'b0011011110010011;
    rom_data[2089]=16'b0010111100000010;
    rom_data[2090]=16'b0011011101011111;
    rom_data[2091]=16'b0010111011101010;
    rom_data[2092]=16'b0011011100101100;
    rom_data[2093]=16'b0010111011100000;
    rom_data[2094]=16'b0011011011111001;
    rom_data[2095]=16'b0010111011100101;
    rom_data[2096]=16'b0011011011000110;
    rom_data[2097]=16'b0010111011111000;
    rom_data[2098]=16'b0011011010010100;
    rom_data[2099]=16'b0010111100011010;
    rom_data[2100]=16'b0011011001100010;
    rom_data[2101]=16'b0010111101001010;
    rom_data[2102]=16'b0011011000110001;
    rom_data[2103]=16'b0010111110000111;
    rom_data[2104]=16'b0011011000000001;
    rom_data[2105]=16'b0010111111010011;
    rom_data[2106]=16'b0011010111010001;
    rom_data[2107]=16'b0011000000101011;
    rom_data[2108]=16'b0011010110100001;
    rom_data[2109]=16'b0011000010010001;
    rom_data[2110]=16'b0011010101110011;
    rom_data[2111]=16'b0011000100000010;
    rom_data[2112]=16'b0011010101000100;
    rom_data[2113]=16'b0011000110000000;
    rom_data[2114]=16'b0011010100010111;
    rom_data[2115]=16'b0011001000001001;
    rom_data[2116]=16'b0011010011101010;
    rom_data[2117]=16'b0011001010011100;
    rom_data[2118]=16'b0011010010111101;
    rom_data[2119]=16'b0011001100111010;
    rom_data[2120]=16'b0011010010010010;
    rom_data[2121]=16'b0011001111100001;
    rom_data[2122]=16'b0011010001100110;
    rom_data[2123]=16'b0011010010010001;
    rom_data[2124]=16'b0011010000111100;
    rom_data[2125]=16'b0011010101001010;
    rom_data[2126]=16'b0011010000010010;
    rom_data[2127]=16'b0011011000001010;
    rom_data[2128]=16'b0011001111101000;
    rom_data[2129]=16'b0011011011010011;
    rom_data[2130]=16'b0011001110111111;
    rom_data[2131]=16'b0011011110100010;
    rom_data[2132]=16'b0011001110010110;
    rom_data[2133]=16'b0011100001111000;
    rom_data[2134]=16'b0011001101101111;
    rom_data[2135]=16'b0011100101010100;
    rom_data[2136]=16'b0011001101000111;
    rom_data[2137]=16'b0011101000110110;
    rom_data[2138]=16'b0011001100100000;
    rom_data[2139]=16'b0011101100011110;
    rom_data[2140]=16'b0011001011111010;
    rom_data[2141]=16'b0011110000001010;
    rom_data[2142]=16'b0011001011010100;
    rom_data[2143]=16'b0011110011111100;
    rom_data[2144]=16'b0011001010101110;
    rom_data[2145]=16'b0011110111110001;
    rom_data[2146]=16'b0011001010001010;
    rom_data[2147]=16'b0011111011101011;
    rom_data[2148]=16'b0011001001100101;
    rom_data[2149]=16'b0011111111101001;
    rom_data[2150]=16'b0011001001000001;
    rom_data[2151]=16'b0100000011101010;
    rom_data[2152]=16'b0011001000011110;
    rom_data[2153]=16'b0100000111101111;
    rom_data[2154]=16'b0011000111111011;
    rom_data[2155]=16'b0100001011110111;
    rom_data[2156]=16'b0011000111011001;
    rom_data[2157]=16'b0100010000000010;
    rom_data[2158]=16'b0011000110110111;
    rom_data[2159]=16'b0100010100001111;
    rom_data[2160]=16'b0011000110010110;
    rom_data[2161]=16'b0100011000100000;
    rom_data[2162]=16'b0011000101110101;
    rom_data[2163]=16'b0100011100110010;
    rom_data[2164]=16'b0011000101010101;
    rom_data[2165]=16'b0100100001000111;
    rom_data[2166]=16'b0011000100110110;
    rom_data[2167]=16'b0100100101011101;
    rom_data[2168]=16'b0011000100010111;
    rom_data[2169]=16'b0100101001110110;
    rom_data[2170]=16'b0011000011111001;
    rom_data[2171]=16'b0100101110010000;
    rom_data[2172]=16'b0011000011011011;
    rom_data[2173]=16'b0100110010101100;
    rom_data[2174]=16'b0011000010111111;
    rom_data[2175]=16'b0100110111001010;
    rom_data[2176]=16'b0011000010100011;
    rom_data[2177]=16'b0100111011101000;
    rom_data[2178]=16'b0011000010001000;
    rom_data[2179]=16'b0101000000001000;
    rom_data[2180]=16'b0011000001101101;
    rom_data[2181]=16'b0101000100101001;
    rom_data[2182]=16'b0011000001010100;
    rom_data[2183]=16'b0101001001001011;
    rom_data[2184]=16'b0011000000111100;
    rom_data[2185]=16'b0101001101101110;
    rom_data[2186]=16'b0011000000100101;
    rom_data[2187]=16'b0101010010010010;
    rom_data[2188]=16'b0011000000001111;
    rom_data[2189]=16'b0101010110110111;
    rom_data[2190]=16'b0010111111111010;
    rom_data[2191]=16'b0101011011011100;
    rom_data[2192]=16'b0010111111111010;
    rom_data[2193]=16'b0101100000000001;
    rom_data[2194]=16'b0011000000001111;
    rom_data[2195]=16'b0101100100100111;
    rom_data[2196]=16'b0011000000100101;
    rom_data[2197]=16'b0101101001001110;
    rom_data[2198]=16'b0011000000111100;
    rom_data[2199]=16'b0101101101110100;
    rom_data[2200]=16'b0011000001010100;
    rom_data[2201]=16'b0101110010011011;

    
// F1
  if (f1_addr==0) begin
    f1_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f1_addr==1) begin
    f1_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f1_addr[0]==1'b0) begin
    f1_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_D_q};
            end

            default: begin
            end
        endcase

   end // if addr=0

// F2
  if (f2_addr==0) begin
    f2_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f2_addr==1) begin
    f2_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f2_addr[0]==1'b0) begin
    f2_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_D_q};
            end

            default: begin
            end
        endcase

   end // if addr=0

// F3
  if (f3_addr==0) begin
    f3_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f3_addr==1) begin
    f3_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f3_addr[0]==1'b0) begin
    f3_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0

// F4
  if (f4_addr==0) begin
    f4_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f4_addr==1) begin
    f4_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f4_addr[0]==1'b0) begin
    f4_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0

// F5
  if (f5_addr==0) begin
    f5_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f5_addr==1) begin
    f5_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f5_addr[0]==1'b0) begin
    f5_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0


// F6
  if (f6_addr==0) begin
    f6_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f6_addr==1) begin
    f6_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f6_addr[0]==1'b0) begin
    f6_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
end // always

always @(posedge f1_addr[0]) begin
    f1_CH_A_q<=f1_CH_A_d;
    f1_CH_B_q<=f1_CH_B_d;
    f1_CH_C_q<=f1_CH_C_d;
    f1_CH_D_q<=f1_CH_D_d;
end

always @(posedge f2_addr[0]) begin
    f2_CH_A_q<=f2_CH_A_d;
    f2_CH_B_q<=f2_CH_B_d;
    f2_CH_C_q<=f2_CH_C_d;
    f2_CH_D_q<=f2_CH_D_d;
end

always @(posedge f3_addr[0]) begin
    f3_CH_A_q<=f3_CH_A_d;
    f3_CH_B_q<=f3_CH_B_d;
    f3_CH_C_q<=f3_CH_C_d;
    f3_CH_D_q<=f3_CH_D_d;
end

always @(posedge f4_addr[0]) begin
    f4_CH_A_q<=f4_CH_A_d;
    f4_CH_B_q<=f4_CH_B_d;
    f4_CH_C_q<=f4_CH_C_d;
    f4_CH_D_q<=f4_CH_D_d;
end

always @(posedge f5_addr[0]) begin
    f5_CH_A_q<=f5_CH_A_d;
    f5_CH_B_q<=f5_CH_B_d;
    f5_CH_C_q<=f5_CH_C_d;
    f5_CH_D_q<=f5_CH_D_d;
end

always @(posedge f6_addr[0]) begin
    f6_CH_A_q<=f6_CH_A_d;
    f6_CH_B_q<=f6_CH_B_d;
    f6_CH_C_q<=f6_CH_C_d;
    f6_CH_D_q<=f6_CH_D_d;
end

always @(posedge clk) begin
    f1_data_q <= f1_data_d;
    f2_data_q <= f2_data_d;
    f3_data_q <= f3_data_d;
    f4_data_q <= f4_data_d;
    f5_data_q <= f5_data_d;
    f6_data_q <= f6_data_d;
end // always
 
endmodule