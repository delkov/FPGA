module mems_rom (
    // INPUT
    input rst,
    input clk,
    input [15:0] f1_addr,
    input [15:0] f2_addr,
    input [15:0] f3_addr,
    input [15:0] f4_addr,
    input [15:0] f5_addr,
    input [15:0] f6_addr,

    input go_home,
    // OUTPUT
    output [23:0] f1_data,
    output [23:0] f2_data,
    output [23:0] f3_data,
    output [23:0] f4_data,
    output [23:0] f5_data,
    output [23:0] f6_data
  );
  
parameter rom_size = 3241;

wire [7:0] rom_data [rom_size:0];


  assign rom_data[ 2]=8'b00101101;
    assign rom_data[ 3]=8'b01011011;
    assign rom_data[ 4]=8'b00101101;
    assign rom_data[ 5]=8'b01011100;
    assign rom_data[ 6]=8'b00101101;
    assign rom_data[ 7]=8'b01011110;
    assign rom_data[ 8]=8'b00101101;
    assign rom_data[ 9]=8'b01011111;
    assign rom_data[10]=8'b00101101;
    assign rom_data[11]=8'b01100001;
    assign rom_data[12]=8'b00101101;
    assign rom_data[13]=8'b01100010;
    assign rom_data[14]=8'b00101101;
    assign rom_data[15]=8'b01100011;
    assign rom_data[16]=8'b00101101;
    assign rom_data[17]=8'b01100101;
    assign rom_data[18]=8'b00101110;
    assign rom_data[19]=8'b01100110;
    assign rom_data[20]=8'b00101110;
    assign rom_data[21]=8'b01100111;
    assign rom_data[22]=8'b00101110;
    assign rom_data[23]=8'b01101001;
    assign rom_data[24]=8'b00101110;
    assign rom_data[25]=8'b01101010;
    assign rom_data[26]=8'b00101110;
    assign rom_data[27]=8'b01101100;
    assign rom_data[28]=8'b00101110;
    assign rom_data[29]=8'b01101101;
    assign rom_data[30]=8'b00101110;
    assign rom_data[31]=8'b01101110;
    assign rom_data[32]=8'b00101110;
    assign rom_data[33]=8'b01110000;
    assign rom_data[34]=8'b00101110;
    assign rom_data[35]=8'b01110001;
    assign rom_data[36]=8'b00101110;
    assign rom_data[37]=8'b01110010;
    assign rom_data[38]=8'b00101110;
    assign rom_data[39]=8'b01110100;
    assign rom_data[40]=8'b00101110;
    assign rom_data[41]=8'b01110101;
    assign rom_data[42]=8'b00101110;
    assign rom_data[43]=8'b01110110;
    assign rom_data[44]=8'b00101110;
    assign rom_data[45]=8'b01110111;
    assign rom_data[46]=8'b00101111;
    assign rom_data[47]=8'b01111001;
    assign rom_data[48]=8'b00101111;
    assign rom_data[49]=8'b01111010;
    assign rom_data[50]=8'b00101111;
    assign rom_data[51]=8'b01111011;
    assign rom_data[52]=8'b00101111;
    assign rom_data[53]=8'b01111100;
    assign rom_data[54]=8'b00101111;
    assign rom_data[55]=8'b01111101;
    assign rom_data[56]=8'b00101111;
    assign rom_data[57]=8'b01111110;
    assign rom_data[58]=8'b00101111;
    assign rom_data[59]=8'b01111111;
    assign rom_data[60]=8'b00101111;
    assign rom_data[61]=8'b10000000;
    assign rom_data[62]=8'b00101111;
    assign rom_data[63]=8'b10000001;
    assign rom_data[64]=8'b00110000;
    assign rom_data[65]=8'b10000010;
    assign rom_data[66]=8'b00110000;
    assign rom_data[67]=8'b10000011;
    assign rom_data[68]=8'b00110000;
    assign rom_data[69]=8'b10000100;
    assign rom_data[70]=8'b00110000;
    assign rom_data[71]=8'b10000101;
    assign rom_data[72]=8'b00110000;
    assign rom_data[73]=8'b10000110;
    assign rom_data[74]=8'b00110000;
    assign rom_data[75]=8'b10000110;
    assign rom_data[76]=8'b00110000;
    assign rom_data[77]=8'b10000111;
    assign rom_data[78]=8'b00110000;
    assign rom_data[79]=8'b10001000;
    assign rom_data[80]=8'b00110000;
    assign rom_data[81]=8'b10001000;
    assign rom_data[82]=8'b00110001;
    assign rom_data[83]=8'b10001001;
    assign rom_data[84]=8'b00110001;
    assign rom_data[85]=8'b10001001;
    assign rom_data[86]=8'b00110001;
    assign rom_data[87]=8'b10001001;
    assign rom_data[88]=8'b00110001;
    assign rom_data[89]=8'b10001010;
    assign rom_data[90]=8'b00110001;
    assign rom_data[91]=8'b10001010;
    assign rom_data[92]=8'b00110001;
    assign rom_data[93]=8'b10001010;
    assign rom_data[94]=8'b00110001;
    assign rom_data[95]=8'b10001010;
    assign rom_data[96]=8'b00110010;
    assign rom_data[97]=8'b10001010;
    assign rom_data[98]=8'b00110010;
    assign rom_data[99]=8'b10001001;
    assign rom_data[100]=8'b00110010;
    assign rom_data[101]=8'b10001001;
    assign rom_data[102]=8'b00110010;
    assign rom_data[103]=8'b10001001;
    assign rom_data[104]=8'b00110010;
    assign rom_data[105]=8'b10001000;
    assign rom_data[106]=8'b00110010;
    assign rom_data[107]=8'b10001000;
    assign rom_data[108]=8'b00110010;
    assign rom_data[109]=8'b10000111;
    assign rom_data[110]=8'b00110010;
    assign rom_data[111]=8'b10000111;
    assign rom_data[112]=8'b00110011;
    assign rom_data[113]=8'b10000110;
    assign rom_data[114]=8'b00110011;
    assign rom_data[115]=8'b10000101;
    assign rom_data[116]=8'b00110011;
    assign rom_data[117]=8'b10000100;
    assign rom_data[118]=8'b00110011;
    assign rom_data[119]=8'b10000011;
    assign rom_data[120]=8'b00110011;
    assign rom_data[121]=8'b10000011;
    assign rom_data[122]=8'b00110011;
    assign rom_data[123]=8'b10000010;
    assign rom_data[124]=8'b00110011;
    assign rom_data[125]=8'b10000001;
    assign rom_data[126]=8'b00110011;
    assign rom_data[127]=8'b10000000;
    assign rom_data[128]=8'b00110100;
    assign rom_data[129]=8'b01111110;
    assign rom_data[130]=8'b00110100;
    assign rom_data[131]=8'b01111101;
    assign rom_data[132]=8'b00110100;
    assign rom_data[133]=8'b01111100;
    assign rom_data[134]=8'b00110100;
    assign rom_data[135]=8'b01111011;
    assign rom_data[136]=8'b00110100;
    assign rom_data[137]=8'b01111010;
    assign rom_data[138]=8'b00110100;
    assign rom_data[139]=8'b01111001;
    assign rom_data[140]=8'b00110100;
    assign rom_data[141]=8'b01110111;
    assign rom_data[142]=8'b00110100;
    assign rom_data[143]=8'b01110110;
    assign rom_data[144]=8'b00110101;
    assign rom_data[145]=8'b01110101;
    assign rom_data[146]=8'b00110101;
    assign rom_data[147]=8'b01110100;
    assign rom_data[148]=8'b00110101;
    assign rom_data[149]=8'b01110010;
    assign rom_data[150]=8'b00110101;
    assign rom_data[151]=8'b01110001;
    assign rom_data[152]=8'b00110101;
    assign rom_data[153]=8'b01110000;
    assign rom_data[154]=8'b00110101;
    assign rom_data[155]=8'b01101110;
    assign rom_data[156]=8'b00110101;
    assign rom_data[157]=8'b01101101;
    assign rom_data[158]=8'b00110101;
    assign rom_data[159]=8'b01101100;
    assign rom_data[160]=8'b00110101;
    assign rom_data[161]=8'b01101010;
    assign rom_data[162]=8'b00110101;
    assign rom_data[163]=8'b01101001;
    assign rom_data[164]=8'b00110110;
    assign rom_data[165]=8'b01101000;
    assign rom_data[166]=8'b00110110;
    assign rom_data[167]=8'b01100110;
    assign rom_data[168]=8'b00110110;
    assign rom_data[169]=8'b01100101;
    assign rom_data[170]=8'b00110110;
    assign rom_data[171]=8'b01100011;
    assign rom_data[172]=8'b00110110;
    assign rom_data[173]=8'b01100010;
    assign rom_data[174]=8'b00110110;
    assign rom_data[175]=8'b01100001;
    assign rom_data[176]=8'b00110110;
    assign rom_data[177]=8'b01011111;
    assign rom_data[178]=8'b00110110;
    assign rom_data[179]=8'b01011110;
    assign rom_data[180]=8'b00110110;
    assign rom_data[181]=8'b01011100;
    assign rom_data[182]=8'b00110110;
    assign rom_data[183]=8'b01011011;
    assign rom_data[184]=8'b00110111;
    assign rom_data[185]=8'b01011010;
    assign rom_data[186]=8'b00110111;
    assign rom_data[187]=8'b01011000;
    assign rom_data[188]=8'b00110111;
    assign rom_data[189]=8'b01010111;
    assign rom_data[190]=8'b00110111;
    assign rom_data[191]=8'b01010101;
    assign rom_data[192]=8'b00110111;
    assign rom_data[193]=8'b01010100;
    assign rom_data[194]=8'b00110111;
    assign rom_data[195]=8'b01010010;
    assign rom_data[196]=8'b00110111;
    assign rom_data[197]=8'b01010001;
    assign rom_data[198]=8'b00110111;
    assign rom_data[199]=8'b01010000;
    assign rom_data[200]=8'b00110111;
    assign rom_data[201]=8'b01001110;
    assign rom_data[202]=8'b00110111;
    assign rom_data[203]=8'b01001101;
    assign rom_data[204]=8'b00111000;
    assign rom_data[205]=8'b01001100;
    assign rom_data[206]=8'b00111000;
    assign rom_data[207]=8'b01001010;
    assign rom_data[208]=8'b00111000;
    assign rom_data[209]=8'b01001001;
    assign rom_data[210]=8'b00111000;
    assign rom_data[211]=8'b01001000;
    assign rom_data[212]=8'b00111000;
    assign rom_data[213]=8'b01000110;
    assign rom_data[214]=8'b00111000;
    assign rom_data[215]=8'b01000101;
    assign rom_data[216]=8'b00111000;
    assign rom_data[217]=8'b01000100;
    assign rom_data[218]=8'b00111000;
    assign rom_data[219]=8'b01000010;
    assign rom_data[220]=8'b00111000;
    assign rom_data[221]=8'b01000001;
    assign rom_data[222]=8'b00111001;
    assign rom_data[223]=8'b01000000;
    assign rom_data[224]=8'b00111001;
    assign rom_data[225]=8'b00111111;
    assign rom_data[226]=8'b00111001;
    assign rom_data[227]=8'b00111101;
    assign rom_data[228]=8'b00111001;
    assign rom_data[229]=8'b00111100;
    assign rom_data[230]=8'b00111001;
    assign rom_data[231]=8'b00111011;
    assign rom_data[232]=8'b00111001;
    assign rom_data[233]=8'b00111010;
    assign rom_data[234]=8'b00111001;
    assign rom_data[235]=8'b00111001;
    assign rom_data[236]=8'b00111001;
    assign rom_data[237]=8'b00111000;
    assign rom_data[238]=8'b00111001;
    assign rom_data[239]=8'b00110110;
    assign rom_data[240]=8'b00111010;
    assign rom_data[241]=8'b00110101;
    assign rom_data[242]=8'b00111010;
    assign rom_data[243]=8'b00110100;
    assign rom_data[244]=8'b00111010;
    assign rom_data[245]=8'b00110011;
    assign rom_data[246]=8'b00111010;
    assign rom_data[247]=8'b00110011;
    assign rom_data[248]=8'b00111010;
    assign rom_data[249]=8'b00110010;
    assign rom_data[250]=8'b00111010;
    assign rom_data[251]=8'b00110001;
    assign rom_data[252]=8'b00111010;
    assign rom_data[253]=8'b00110000;
    assign rom_data[254]=8'b00111010;
    assign rom_data[255]=8'b00101111;
    assign rom_data[256]=8'b00111011;
    assign rom_data[257]=8'b00101111;
    assign rom_data[258]=8'b00111011;
    assign rom_data[259]=8'b00101110;
    assign rom_data[260]=8'b00111011;
    assign rom_data[261]=8'b00101110;
    assign rom_data[262]=8'b00111011;
    assign rom_data[263]=8'b00101101;
    assign rom_data[264]=8'b00111011;
    assign rom_data[265]=8'b00101101;
    assign rom_data[266]=8'b00111011;
    assign rom_data[267]=8'b00101100;
    assign rom_data[268]=8'b00111011;
    assign rom_data[269]=8'b00101100;
    assign rom_data[270]=8'b00111100;
    assign rom_data[271]=8'b00101100;
    assign rom_data[272]=8'b00111100;
    assign rom_data[273]=8'b00101100;
    assign rom_data[274]=8'b00111100;
    assign rom_data[275]=8'b00101100;
    assign rom_data[276]=8'b00111100;
    assign rom_data[277]=8'b00101100;
    assign rom_data[278]=8'b00111100;
    assign rom_data[279]=8'b00101100;
    assign rom_data[280]=8'b00111100;
    assign rom_data[281]=8'b00101101;
    assign rom_data[282]=8'b00111100;
    assign rom_data[283]=8'b00101101;
    assign rom_data[284]=8'b00111100;
    assign rom_data[285]=8'b00101101;
    assign rom_data[286]=8'b00111101;
    assign rom_data[287]=8'b00101110;
    assign rom_data[288]=8'b00111101;
    assign rom_data[289]=8'b00101111;
    assign rom_data[290]=8'b00111101;
    assign rom_data[291]=8'b00101111;
    assign rom_data[292]=8'b00111101;
    assign rom_data[293]=8'b00110000;
    assign rom_data[294]=8'b00111101;
    assign rom_data[295]=8'b00110001;
    assign rom_data[296]=8'b00111101;
    assign rom_data[297]=8'b00110001;
    assign rom_data[298]=8'b00111101;
    assign rom_data[299]=8'b00110010;
    assign rom_data[300]=8'b00111110;
    assign rom_data[301]=8'b00110011;
    assign rom_data[302]=8'b00111110;
    assign rom_data[303]=8'b00110100;
    assign rom_data[304]=8'b00111110;
    assign rom_data[305]=8'b00110101;
    assign rom_data[306]=8'b00111110;
    assign rom_data[307]=8'b00110110;
    assign rom_data[308]=8'b00111110;
    assign rom_data[309]=8'b00110111;
    assign rom_data[310]=8'b00111110;
    assign rom_data[311]=8'b00111000;
    assign rom_data[312]=8'b00111110;
    assign rom_data[313]=8'b00111010;
    assign rom_data[314]=8'b00111110;
    assign rom_data[315]=8'b00111011;
    assign rom_data[316]=8'b00111110;
    assign rom_data[317]=8'b00111100;
    assign rom_data[318]=8'b00111111;
    assign rom_data[319]=8'b00111101;
    assign rom_data[320]=8'b00111111;
    assign rom_data[321]=8'b00111110;
    assign rom_data[322]=8'b00111111;
    assign rom_data[323]=8'b01000000;
    assign rom_data[324]=8'b00111111;
    assign rom_data[325]=8'b01000001;
    assign rom_data[326]=8'b00111111;
    assign rom_data[327]=8'b01000010;
    assign rom_data[328]=8'b00111111;
    assign rom_data[329]=8'b01000100;
    assign rom_data[330]=8'b00111111;
    assign rom_data[331]=8'b01000101;
    assign rom_data[332]=8'b00111111;
    assign rom_data[333]=8'b01000110;
    assign rom_data[334]=8'b00111111;
    assign rom_data[335]=8'b01000111;
    assign rom_data[336]=8'b01000000;
    assign rom_data[337]=8'b01001001;
    assign rom_data[338]=8'b01000000;
    assign rom_data[339]=8'b01001010;
    assign rom_data[340]=8'b01000000;
    assign rom_data[341]=8'b01001100;
    assign rom_data[342]=8'b01000000;
    assign rom_data[343]=8'b01001101;
    assign rom_data[344]=8'b01000000;
    assign rom_data[345]=8'b01001110;
    assign rom_data[346]=8'b01000000;
    assign rom_data[347]=8'b01010000;
    assign rom_data[348]=8'b01000000;
    assign rom_data[349]=8'b01010001;
    assign rom_data[350]=8'b01000000;
    assign rom_data[351]=8'b01010010;
    assign rom_data[352]=8'b01000000;
    assign rom_data[353]=8'b01010100;
    assign rom_data[354]=8'b01000000;
    assign rom_data[355]=8'b01010101;
    assign rom_data[356]=8'b01000001;
    assign rom_data[357]=8'b01010111;
    assign rom_data[358]=8'b01000001;
    assign rom_data[359]=8'b01011000;
    assign rom_data[360]=8'b01000001;
    assign rom_data[361]=8'b01011010;
    assign rom_data[362]=8'b01000001;
    assign rom_data[363]=8'b01011011;
    assign rom_data[364]=8'b01000001;
    assign rom_data[365]=8'b01011100;
    assign rom_data[366]=8'b01000001;
    assign rom_data[367]=8'b01011110;
    assign rom_data[368]=8'b01000001;
    assign rom_data[369]=8'b01011111;
    assign rom_data[370]=8'b01000001;
    assign rom_data[371]=8'b01100001;
    assign rom_data[372]=8'b01000001;
    assign rom_data[373]=8'b01100010;
    assign rom_data[374]=8'b01000001;
    assign rom_data[375]=8'b01100011;
    assign rom_data[376]=8'b01000010;
    assign rom_data[377]=8'b01100101;
    assign rom_data[378]=8'b01000010;
    assign rom_data[379]=8'b01100110;
    assign rom_data[380]=8'b01000010;
    assign rom_data[381]=8'b01100111;
    assign rom_data[382]=8'b01000010;
    assign rom_data[383]=8'b01101001;
    assign rom_data[384]=8'b01000010;
    assign rom_data[385]=8'b01101010;
    assign rom_data[386]=8'b01000010;
    assign rom_data[387]=8'b01101100;
    assign rom_data[388]=8'b01000010;
    assign rom_data[389]=8'b01101101;
    assign rom_data[390]=8'b01000010;
    assign rom_data[391]=8'b01101110;
    assign rom_data[392]=8'b01000010;
    assign rom_data[393]=8'b01110000;
    assign rom_data[394]=8'b01000011;
    assign rom_data[395]=8'b01110001;
    assign rom_data[396]=8'b01000011;
    assign rom_data[397]=8'b01110010;
    assign rom_data[398]=8'b01000011;
    assign rom_data[399]=8'b01110100;
    assign rom_data[400]=8'b01000011;
    assign rom_data[401]=8'b01110101;
    assign rom_data[402]=8'b01000011;
    assign rom_data[403]=8'b01110110;
    assign rom_data[404]=8'b01000011;
    assign rom_data[405]=8'b01110111;
    assign rom_data[406]=8'b01000011;
    assign rom_data[407]=8'b01111001;
    assign rom_data[408]=8'b01000011;
    assign rom_data[409]=8'b01111010;
    assign rom_data[410]=8'b01000011;
    assign rom_data[411]=8'b01111011;
    assign rom_data[412]=8'b01000011;
    assign rom_data[413]=8'b01111100;
    assign rom_data[414]=8'b01000100;
    assign rom_data[415]=8'b01111101;
    assign rom_data[416]=8'b01000100;
    assign rom_data[417]=8'b01111110;
    assign rom_data[418]=8'b01000100;
    assign rom_data[419]=8'b01111111;
    assign rom_data[420]=8'b01000100;
    assign rom_data[421]=8'b10000000;
    assign rom_data[422]=8'b01000100;
    assign rom_data[423]=8'b10000001;
    assign rom_data[424]=8'b01000100;
    assign rom_data[425]=8'b10000010;
    assign rom_data[426]=8'b01000100;
    assign rom_data[427]=8'b10000011;
    assign rom_data[428]=8'b01000100;
    assign rom_data[429]=8'b10000100;
    assign rom_data[430]=8'b01000101;
    assign rom_data[431]=8'b10000101;
    assign rom_data[432]=8'b01000101;
    assign rom_data[433]=8'b10000110;
    assign rom_data[434]=8'b01000101;
    assign rom_data[435]=8'b10000110;
    assign rom_data[436]=8'b01000101;
    assign rom_data[437]=8'b10000111;
    assign rom_data[438]=8'b01000101;
    assign rom_data[439]=8'b10001000;
    assign rom_data[440]=8'b01000101;
    assign rom_data[441]=8'b10001000;
    assign rom_data[442]=8'b01000101;
    assign rom_data[443]=8'b10001001;
    assign rom_data[444]=8'b01000110;
    assign rom_data[445]=8'b10001001;
    assign rom_data[446]=8'b01000110;
    assign rom_data[447]=8'b10001001;
    assign rom_data[448]=8'b01000110;
    assign rom_data[449]=8'b10001010;
    assign rom_data[450]=8'b01000110;
    assign rom_data[451]=8'b10001010;
    assign rom_data[452]=8'b01000110;
    assign rom_data[453]=8'b10001010;
    assign rom_data[454]=8'b01000110;
    assign rom_data[455]=8'b10001010;
    assign rom_data[456]=8'b01000110;
    assign rom_data[457]=8'b10001010;
    assign rom_data[458]=8'b01000111;
    assign rom_data[459]=8'b10001001;
    assign rom_data[460]=8'b01000111;
    assign rom_data[461]=8'b10001001;
    assign rom_data[462]=8'b01000111;
    assign rom_data[463]=8'b10001001;
    assign rom_data[464]=8'b01000111;
    assign rom_data[465]=8'b10001000;
    assign rom_data[466]=8'b01000111;
    assign rom_data[467]=8'b10001000;
    assign rom_data[468]=8'b01000111;
    assign rom_data[469]=8'b10000111;
    assign rom_data[470]=8'b01000111;
    assign rom_data[471]=8'b10000111;
    assign rom_data[472]=8'b01000111;
    assign rom_data[473]=8'b10000110;
    assign rom_data[474]=8'b01001000;
    assign rom_data[475]=8'b10000101;
    assign rom_data[476]=8'b01001000;
    assign rom_data[477]=8'b10000100;
    assign rom_data[478]=8'b01001000;
    assign rom_data[479]=8'b10000011;
    assign rom_data[480]=8'b01001000;
    assign rom_data[481]=8'b10000011;
    assign rom_data[482]=8'b01001000;
    assign rom_data[483]=8'b10000010;
    assign rom_data[484]=8'b01001000;
    assign rom_data[485]=8'b10000001;
    assign rom_data[486]=8'b01001000;
    assign rom_data[487]=8'b10000000;
    assign rom_data[488]=8'b01001000;
    assign rom_data[489]=8'b01111110;
    assign rom_data[490]=8'b01001001;
    assign rom_data[491]=8'b01111101;
    assign rom_data[492]=8'b01001001;
    assign rom_data[493]=8'b01111100;
    assign rom_data[494]=8'b01001001;
    assign rom_data[495]=8'b01111011;
    assign rom_data[496]=8'b01001001;
    assign rom_data[497]=8'b01111010;
    assign rom_data[498]=8'b01001001;
    assign rom_data[499]=8'b01111001;
    assign rom_data[500]=8'b01001001;
    assign rom_data[501]=8'b01110111;
    assign rom_data[502]=8'b01001001;
    assign rom_data[503]=8'b01110110;
    assign rom_data[504]=8'b01001001;
    assign rom_data[505]=8'b01110101;
    assign rom_data[506]=8'b01001001;
    assign rom_data[507]=8'b01110100;
    assign rom_data[508]=8'b01001010;
    assign rom_data[509]=8'b01110010;
    assign rom_data[510]=8'b01001010;
    assign rom_data[511]=8'b01110001;
    assign rom_data[512]=8'b01001010;
    assign rom_data[513]=8'b01110000;
    assign rom_data[514]=8'b01001010;
    assign rom_data[515]=8'b01101110;
    assign rom_data[516]=8'b01001010;
    assign rom_data[517]=8'b01101101;
    assign rom_data[518]=8'b01001010;
    assign rom_data[519]=8'b01101100;
    assign rom_data[520]=8'b01001010;
    assign rom_data[521]=8'b01101010;
    assign rom_data[522]=8'b01001010;
    assign rom_data[523]=8'b01101001;
    assign rom_data[524]=8'b01001010;
    assign rom_data[525]=8'b01101000;
    assign rom_data[526]=8'b01001011;
    assign rom_data[527]=8'b01100110;
    assign rom_data[528]=8'b01001011;
    assign rom_data[529]=8'b01100101;
    assign rom_data[530]=8'b01001011;
    assign rom_data[531]=8'b01100011;
    assign rom_data[532]=8'b01001011;
    assign rom_data[533]=8'b01100010;
    assign rom_data[534]=8'b01001011;
    assign rom_data[535]=8'b01100001;
    assign rom_data[536]=8'b01001011;
    assign rom_data[537]=8'b01011111;
    assign rom_data[538]=8'b01001011;
    assign rom_data[539]=8'b01011110;
    assign rom_data[540]=8'b01001011;
    assign rom_data[541]=8'b01011100;
    assign rom_data[542]=8'b01001011;
    assign rom_data[543]=8'b01011011;
    assign rom_data[544]=8'b01001011;
    assign rom_data[545]=8'b01011001;
    assign rom_data[546]=8'b01001100;
    assign rom_data[547]=8'b01011000;
    assign rom_data[548]=8'b01001100;
    assign rom_data[549]=8'b01010111;
    assign rom_data[550]=8'b01001100;
    assign rom_data[551]=8'b01010101;
    assign rom_data[552]=8'b01001100;
    assign rom_data[553]=8'b01010100;
    assign rom_data[554]=8'b01001100;
    assign rom_data[555]=8'b01010010;
    assign rom_data[556]=8'b01001100;
    assign rom_data[557]=8'b01010001;
    assign rom_data[558]=8'b01001100;
    assign rom_data[559]=8'b01010000;
    assign rom_data[560]=8'b01001100;
    assign rom_data[561]=8'b01001110;
    assign rom_data[562]=8'b01001100;
    assign rom_data[563]=8'b01001101;
    assign rom_data[564]=8'b01001100;
    assign rom_data[565]=8'b01001100;
    assign rom_data[566]=8'b01001101;
    assign rom_data[567]=8'b01001010;
    assign rom_data[568]=8'b01001101;
    assign rom_data[569]=8'b01001001;
    assign rom_data[570]=8'b01001101;
    assign rom_data[571]=8'b01001000;
    assign rom_data[572]=8'b01001101;
    assign rom_data[573]=8'b01000110;
    assign rom_data[574]=8'b01001101;
    assign rom_data[575]=8'b01000101;
    assign rom_data[576]=8'b01001101;
    assign rom_data[577]=8'b01000100;
    assign rom_data[578]=8'b01001101;
    assign rom_data[579]=8'b01000010;
    assign rom_data[580]=8'b01001101;
    assign rom_data[581]=8'b01000001;
    assign rom_data[582]=8'b01001101;
    assign rom_data[583]=8'b01000000;
    assign rom_data[584]=8'b01001101;
    assign rom_data[585]=8'b00111111;
    assign rom_data[586]=8'b01001110;
    assign rom_data[587]=8'b00111101;
    assign rom_data[588]=8'b01001110;
    assign rom_data[589]=8'b00111100;
    assign rom_data[590]=8'b01001110;
    assign rom_data[591]=8'b00111011;
    assign rom_data[592]=8'b01001110;
    assign rom_data[593]=8'b00111010;
    assign rom_data[594]=8'b01001110;
    assign rom_data[595]=8'b00111001;
    assign rom_data[596]=8'b01001110;
    assign rom_data[597]=8'b00111000;
    assign rom_data[598]=8'b01001110;
    assign rom_data[599]=8'b00110110;
    assign rom_data[600]=8'b01001110;
    assign rom_data[601]=8'b00110101;
    assign rom_data[602]=8'b01001111;
    assign rom_data[603]=8'b00110100;
    assign rom_data[604]=8'b01001111;
    assign rom_data[605]=8'b00110011;
    assign rom_data[606]=8'b01001111;
    assign rom_data[607]=8'b00110011;
    assign rom_data[608]=8'b01001111;
    assign rom_data[609]=8'b00110010;
    assign rom_data[610]=8'b01001111;
    assign rom_data[611]=8'b00110001;
    assign rom_data[612]=8'b01001111;
    assign rom_data[613]=8'b00110000;
    assign rom_data[614]=8'b01001111;
    assign rom_data[615]=8'b00101111;
    assign rom_data[616]=8'b01001111;
    assign rom_data[617]=8'b00101111;
    assign rom_data[618]=8'b01010000;
    assign rom_data[619]=8'b00101110;
    assign rom_data[620]=8'b01010000;
    assign rom_data[621]=8'b00101110;
    assign rom_data[622]=8'b01010000;
    assign rom_data[623]=8'b00101101;
    assign rom_data[624]=8'b01010000;
    assign rom_data[625]=8'b00101101;
    assign rom_data[626]=8'b01010000;
    assign rom_data[627]=8'b00101100;
    assign rom_data[628]=8'b01010000;
    assign rom_data[629]=8'b00101100;
    assign rom_data[630]=8'b01010000;
    assign rom_data[631]=8'b00101100;
    assign rom_data[632]=8'b01010001;
    assign rom_data[633]=8'b00101100;
    assign rom_data[634]=8'b01010001;
    assign rom_data[635]=8'b00101100;
    assign rom_data[636]=8'b01010001;
    assign rom_data[637]=8'b00101100;
    assign rom_data[638]=8'b01010001;
    assign rom_data[639]=8'b00101100;
    assign rom_data[640]=8'b01010001;
    assign rom_data[641]=8'b00101101;
    assign rom_data[642]=8'b01010001;
    assign rom_data[643]=8'b00101101;
    assign rom_data[644]=8'b01010001;
    assign rom_data[645]=8'b00101101;
    assign rom_data[646]=8'b01010001;
    assign rom_data[647]=8'b00101110;
    assign rom_data[648]=8'b01010010;
    assign rom_data[649]=8'b00101111;
    assign rom_data[650]=8'b01010010;
    assign rom_data[651]=8'b00101111;
    assign rom_data[652]=8'b01010010;
    assign rom_data[653]=8'b00110000;
    assign rom_data[654]=8'b01010010;
    assign rom_data[655]=8'b00110001;
    assign rom_data[656]=8'b01010010;
    assign rom_data[657]=8'b00110001;
    assign rom_data[658]=8'b01010010;
    assign rom_data[659]=8'b00110010;
    assign rom_data[660]=8'b01010010;
    assign rom_data[661]=8'b00110011;
    assign rom_data[662]=8'b01010011;
    assign rom_data[663]=8'b00110100;
    assign rom_data[664]=8'b01010011;
    assign rom_data[665]=8'b00110101;
    assign rom_data[666]=8'b01010011;
    assign rom_data[667]=8'b00110110;
    assign rom_data[668]=8'b01010011;
    assign rom_data[669]=8'b00110111;
    assign rom_data[670]=8'b01010011;
    assign rom_data[671]=8'b00111000;
    assign rom_data[672]=8'b01010011;
    assign rom_data[673]=8'b00111010;
    assign rom_data[674]=8'b01010011;
    assign rom_data[675]=8'b00111011;
    assign rom_data[676]=8'b01010011;
    assign rom_data[677]=8'b00111100;
    assign rom_data[678]=8'b01010011;
    assign rom_data[679]=8'b00111101;
    assign rom_data[680]=8'b01010100;
    assign rom_data[681]=8'b00111110;
    assign rom_data[682]=8'b01010100;
    assign rom_data[683]=8'b01000000;
    assign rom_data[684]=8'b01010100;
    assign rom_data[685]=8'b01000001;
    assign rom_data[686]=8'b01010100;
    assign rom_data[687]=8'b01000010;
    assign rom_data[688]=8'b01010100;
    assign rom_data[689]=8'b01000100;
    assign rom_data[690]=8'b01010100;
    assign rom_data[691]=8'b01000101;
    assign rom_data[692]=8'b01010100;
    assign rom_data[693]=8'b01000110;
    assign rom_data[694]=8'b01010100;
    assign rom_data[695]=8'b01000111;
    assign rom_data[696]=8'b01010100;
    assign rom_data[697]=8'b01001001;
    assign rom_data[698]=8'b01010101;
    assign rom_data[699]=8'b01001010;
    assign rom_data[700]=8'b01010101;
    assign rom_data[701]=8'b01001100;
    assign rom_data[702]=8'b01010101;
    assign rom_data[703]=8'b01001101;
    assign rom_data[704]=8'b01010101;
    assign rom_data[705]=8'b01001110;
    assign rom_data[706]=8'b01010101;
    assign rom_data[707]=8'b01010000;
    assign rom_data[708]=8'b01010101;
    assign rom_data[709]=8'b01010001;
    assign rom_data[710]=8'b01010101;
    assign rom_data[711]=8'b01010010;
    assign rom_data[712]=8'b01010101;
    assign rom_data[713]=8'b01010100;
    assign rom_data[714]=8'b01010101;
    assign rom_data[715]=8'b01010101;
    assign rom_data[716]=8'b01010101;
    assign rom_data[717]=8'b01010111;
    assign rom_data[718]=8'b01010110;
    assign rom_data[719]=8'b01011000;
    assign rom_data[720]=8'b01010110;
    assign rom_data[721]=8'b01011010;
    assign rom_data[722]=8'b01010110;
    assign rom_data[723]=8'b01011011;
    assign rom_data[724]=8'b01010110;
    assign rom_data[725]=8'b01011100;
    assign rom_data[726]=8'b01010110;
    assign rom_data[727]=8'b01011110;
    assign rom_data[728]=8'b01010110;
    assign rom_data[729]=8'b01011111;
    assign rom_data[730]=8'b01010110;
    assign rom_data[731]=8'b01100001;
    assign rom_data[732]=8'b01010110;
    assign rom_data[733]=8'b01100010;
    assign rom_data[734]=8'b01010110;
    assign rom_data[735]=8'b01100011;
    assign rom_data[736]=8'b01010110;
    assign rom_data[737]=8'b01100101;
    assign rom_data[738]=8'b01010111;
    assign rom_data[739]=8'b01100110;
    assign rom_data[740]=8'b01010111;
    assign rom_data[741]=8'b01100111;
    assign rom_data[742]=8'b01010111;
    assign rom_data[743]=8'b01101001;
    assign rom_data[744]=8'b01010111;
    assign rom_data[745]=8'b01101010;
    assign rom_data[746]=8'b01010111;
    assign rom_data[747]=8'b01101100;
    assign rom_data[748]=8'b01010111;
    assign rom_data[749]=8'b01101101;
    assign rom_data[750]=8'b01010111;
    assign rom_data[751]=8'b01101110;
    assign rom_data[752]=8'b01010111;
    assign rom_data[753]=8'b01110000;
    assign rom_data[754]=8'b01010111;
    assign rom_data[755]=8'b01110001;
    assign rom_data[756]=8'b01010111;
    assign rom_data[757]=8'b01110010;
    assign rom_data[758]=8'b01011000;
    assign rom_data[759]=8'b01110100;
    assign rom_data[760]=8'b01011000;
    assign rom_data[761]=8'b01110101;
    assign rom_data[762]=8'b01011000;
    assign rom_data[763]=8'b01110110;
    assign rom_data[764]=8'b01011000;
    assign rom_data[765]=8'b01110111;
    assign rom_data[766]=8'b01011000;
    assign rom_data[767]=8'b01111001;
    assign rom_data[768]=8'b01011000;
    assign rom_data[769]=8'b01111010;
    assign rom_data[770]=8'b01011000;
    assign rom_data[771]=8'b01111011;
    assign rom_data[772]=8'b01011000;
    assign rom_data[773]=8'b01111100;
    assign rom_data[774]=8'b01011000;
    assign rom_data[775]=8'b01111101;
    assign rom_data[776]=8'b01011001;
    assign rom_data[777]=8'b01111110;
    assign rom_data[778]=8'b01011001;
    assign rom_data[779]=8'b01111111;
    assign rom_data[780]=8'b01011001;
    assign rom_data[781]=8'b10000000;
    assign rom_data[782]=8'b01011001;
    assign rom_data[783]=8'b10000001;
    assign rom_data[784]=8'b01011001;
    assign rom_data[785]=8'b10000010;
    assign rom_data[786]=8'b01011001;
    assign rom_data[787]=8'b10000011;
    assign rom_data[788]=8'b01011001;
    assign rom_data[789]=8'b10000100;
    assign rom_data[790]=8'b01011001;
    assign rom_data[791]=8'b10000101;
    assign rom_data[792]=8'b01011010;
    assign rom_data[793]=8'b10000110;
    assign rom_data[794]=8'b01011010;
    assign rom_data[795]=8'b10000110;
    assign rom_data[796]=8'b01011010;
    assign rom_data[797]=8'b10000111;
    assign rom_data[798]=8'b01011010;
    assign rom_data[799]=8'b10001000;
    assign rom_data[800]=8'b01011010;
    assign rom_data[801]=8'b10001000;
    assign rom_data[802]=8'b01011010;
    assign rom_data[803]=8'b10001001;
    assign rom_data[804]=8'b01011010;
    assign rom_data[805]=8'b10001001;
    assign rom_data[806]=8'b01011011;
    assign rom_data[807]=8'b10001001;
    assign rom_data[808]=8'b01011011;
    assign rom_data[809]=8'b10001010;
    assign rom_data[810]=8'b01011011;
    assign rom_data[811]=8'b10001010;
    assign rom_data[812]=8'b01011011;
    assign rom_data[813]=8'b10001010;
    assign rom_data[814]=8'b01011011;
    assign rom_data[815]=8'b10001010;
    assign rom_data[816]=8'b01011011;
    assign rom_data[817]=8'b10001010;
    assign rom_data[818]=8'b01011011;
    assign rom_data[819]=8'b10001001;
    assign rom_data[820]=8'b01011011;
    assign rom_data[821]=8'b10001001;
    assign rom_data[822]=8'b01011100;
    assign rom_data[823]=8'b10001001;
    assign rom_data[824]=8'b01011100;
    assign rom_data[825]=8'b10001000;
    assign rom_data[826]=8'b01011100;
    assign rom_data[827]=8'b10001000;
    assign rom_data[828]=8'b01011100;
    assign rom_data[829]=8'b10000111;
    assign rom_data[830]=8'b01011100;
    assign rom_data[831]=8'b10000111;
    assign rom_data[832]=8'b01011100;
    assign rom_data[833]=8'b10000110;
    assign rom_data[834]=8'b01011100;
    assign rom_data[835]=8'b10000101;
    assign rom_data[836]=8'b01011101;
    assign rom_data[837]=8'b10000100;
    assign rom_data[838]=8'b01011101;
    assign rom_data[839]=8'b10000011;
    assign rom_data[840]=8'b01011101;
    assign rom_data[841]=8'b10000011;
    assign rom_data[842]=8'b01011101;
    assign rom_data[843]=8'b10000010;
    assign rom_data[844]=8'b01011101;
    assign rom_data[845]=8'b10000001;
    assign rom_data[846]=8'b01011101;
    assign rom_data[847]=8'b10000000;
    assign rom_data[848]=8'b01011101;
    assign rom_data[849]=8'b01111110;
    assign rom_data[850]=8'b01011101;
    assign rom_data[851]=8'b01111101;
    assign rom_data[852]=8'b01011110;
    assign rom_data[853]=8'b01111100;
    assign rom_data[854]=8'b01011110;
    assign rom_data[855]=8'b01111011;
    assign rom_data[856]=8'b01011110;
    assign rom_data[857]=8'b01111010;
    assign rom_data[858]=8'b01011110;
    assign rom_data[859]=8'b01111001;
    assign rom_data[860]=8'b01011110;
    assign rom_data[861]=8'b01110111;
    assign rom_data[862]=8'b01011110;
    assign rom_data[863]=8'b01110110;
    assign rom_data[864]=8'b01011110;
    assign rom_data[865]=8'b01110101;
    assign rom_data[866]=8'b01011110;
    assign rom_data[867]=8'b01110100;
    assign rom_data[868]=8'b01011110;
    assign rom_data[869]=8'b01110010;
    assign rom_data[870]=8'b01011111;
    assign rom_data[871]=8'b01110001;
    assign rom_data[872]=8'b01011111;
    assign rom_data[873]=8'b01110000;
    assign rom_data[874]=8'b01011111;
    assign rom_data[875]=8'b01101110;
    assign rom_data[876]=8'b01011111;
    assign rom_data[877]=8'b01101101;
    assign rom_data[878]=8'b01011111;
    assign rom_data[879]=8'b01101100;
    assign rom_data[880]=8'b01011111;
    assign rom_data[881]=8'b01101010;
    assign rom_data[882]=8'b01011111;
    assign rom_data[883]=8'b01101001;
    assign rom_data[884]=8'b01011111;
    assign rom_data[885]=8'b01101000;
    assign rom_data[886]=8'b01011111;
    assign rom_data[887]=8'b01100110;
    assign rom_data[888]=8'b01011111;
    assign rom_data[889]=8'b01100101;
    assign rom_data[890]=8'b01100000;
    assign rom_data[891]=8'b01100011;
    assign rom_data[892]=8'b01100000;
    assign rom_data[893]=8'b01100010;
    assign rom_data[894]=8'b01100000;
    assign rom_data[895]=8'b01100001;
    assign rom_data[896]=8'b01100000;
    assign rom_data[897]=8'b01011111;
    assign rom_data[898]=8'b01100000;
    assign rom_data[899]=8'b01011110;
    assign rom_data[900]=8'b01100000;
    assign rom_data[901]=8'b01011100;
    assign rom_data[902]=8'b01100000;
    assign rom_data[903]=8'b01011011;
    assign rom_data[904]=8'b01100000;
    assign rom_data[905]=8'b01011001;
    assign rom_data[906]=8'b01100000;
    assign rom_data[907]=8'b01011000;
    assign rom_data[908]=8'b01100000;
    assign rom_data[909]=8'b01010111;
    assign rom_data[910]=8'b01100001;
    assign rom_data[911]=8'b01010101;
    assign rom_data[912]=8'b01100001;
    assign rom_data[913]=8'b01010100;
    assign rom_data[914]=8'b01100001;
    assign rom_data[915]=8'b01010010;
    assign rom_data[916]=8'b01100001;
    assign rom_data[917]=8'b01010001;
    assign rom_data[918]=8'b01100001;
    assign rom_data[919]=8'b01010000;
    assign rom_data[920]=8'b01100001;
    assign rom_data[921]=8'b01001110;
    assign rom_data[922]=8'b01100001;
    assign rom_data[923]=8'b01001101;
    assign rom_data[924]=8'b01100001;
    assign rom_data[925]=8'b01001100;
    assign rom_data[926]=8'b01100001;
    assign rom_data[927]=8'b01001010;
    assign rom_data[928]=8'b01100001;
    assign rom_data[929]=8'b01001001;
    assign rom_data[930]=8'b01100010;
    assign rom_data[931]=8'b01001000;
    assign rom_data[932]=8'b01100010;
    assign rom_data[933]=8'b01000110;
    assign rom_data[934]=8'b01100010;
    assign rom_data[935]=8'b01000101;
    assign rom_data[936]=8'b01100010;
    assign rom_data[937]=8'b01000100;
    assign rom_data[938]=8'b01100010;
    assign rom_data[939]=8'b01000010;
    assign rom_data[940]=8'b01100010;
    assign rom_data[941]=8'b01000001;
    assign rom_data[942]=8'b01100010;
    assign rom_data[943]=8'b01000000;
    assign rom_data[944]=8'b01100010;
    assign rom_data[945]=8'b00111111;
    assign rom_data[946]=8'b01100010;
    assign rom_data[947]=8'b00111101;
    assign rom_data[948]=8'b01100011;
    assign rom_data[949]=8'b00111100;
    assign rom_data[950]=8'b01100011;
    assign rom_data[951]=8'b00111011;
    assign rom_data[952]=8'b01100011;
    assign rom_data[953]=8'b00111010;
    assign rom_data[954]=8'b01100011;
    assign rom_data[955]=8'b00111001;
    assign rom_data[956]=8'b01100011;
    assign rom_data[957]=8'b00111000;
    assign rom_data[958]=8'b01100011;
    assign rom_data[959]=8'b00110110;
    assign rom_data[960]=8'b01100011;
    assign rom_data[961]=8'b00110101;
    assign rom_data[962]=8'b01100011;
    assign rom_data[963]=8'b00110100;
    assign rom_data[964]=8'b01100011;
    assign rom_data[965]=8'b00110011;
    assign rom_data[966]=8'b01100100;
    assign rom_data[967]=8'b00110011;
    assign rom_data[968]=8'b01100100;
    assign rom_data[969]=8'b00110010;
    assign rom_data[970]=8'b01100100;
    assign rom_data[971]=8'b00110001;
    assign rom_data[972]=8'b01100100;
    assign rom_data[973]=8'b00110000;
    assign rom_data[974]=8'b01100100;
    assign rom_data[975]=8'b00101111;
    assign rom_data[976]=8'b01100100;
    assign rom_data[977]=8'b00101111;
    assign rom_data[978]=8'b01100100;
    assign rom_data[979]=8'b00101110;
    assign rom_data[980]=8'b01100101;
    assign rom_data[981]=8'b00101110;
    assign rom_data[982]=8'b01100101;
    assign rom_data[983]=8'b00101101;
    assign rom_data[984]=8'b01100101;
    assign rom_data[985]=8'b00101101;
    assign rom_data[986]=8'b01100101;
    assign rom_data[987]=8'b00101100;
    assign rom_data[988]=8'b01100101;
    assign rom_data[989]=8'b00101100;
    assign rom_data[990]=8'b01100101;
    assign rom_data[991]=8'b00101100;
    assign rom_data[992]=8'b01100101;
    assign rom_data[993]=8'b00101100;
    assign rom_data[994]=8'b01100110;
    assign rom_data[995]=8'b00101100;
    assign rom_data[996]=8'b01100110;
    assign rom_data[997]=8'b00101100;
    assign rom_data[998]=8'b01100110;
    assign rom_data[999]=8'b00101100;
    assign rom_data[1000]=8'b01100110;
    assign rom_data[1001]=8'b00101101;
    assign rom_data[1002]=8'b01100110;
    assign rom_data[1003]=8'b00101101;
    assign rom_data[1004]=8'b01100110;
    assign rom_data[1005]=8'b00101101;
    assign rom_data[1006]=8'b01100110;
    assign rom_data[1007]=8'b00101110;
    assign rom_data[1008]=8'b01100110;
    assign rom_data[1009]=8'b00101111;
    assign rom_data[1010]=8'b01100111;
    assign rom_data[1011]=8'b00101111;
    assign rom_data[1012]=8'b01100111;
    assign rom_data[1013]=8'b00110000;
    assign rom_data[1014]=8'b01100111;
    assign rom_data[1015]=8'b00110001;
    assign rom_data[1016]=8'b01100111;
    assign rom_data[1017]=8'b00110001;
    assign rom_data[1018]=8'b01100111;
    assign rom_data[1019]=8'b00110010;
    assign rom_data[1020]=8'b01100111;
    assign rom_data[1021]=8'b00110011;
    assign rom_data[1022]=8'b01100111;
    assign rom_data[1023]=8'b00110100;
    assign rom_data[1024]=8'b01101000;
    assign rom_data[1025]=8'b00110101;
    assign rom_data[1026]=8'b01101000;
    assign rom_data[1027]=8'b00110110;
    assign rom_data[1028]=8'b01101000;
    assign rom_data[1029]=8'b00110111;
    assign rom_data[1030]=8'b01101000;
    assign rom_data[1031]=8'b00111000;
    assign rom_data[1032]=8'b01101000;
    assign rom_data[1033]=8'b00111010;
    assign rom_data[1034]=8'b01101000;
    assign rom_data[1035]=8'b00111011;
    assign rom_data[1036]=8'b01101000;
    assign rom_data[1037]=8'b00111100;
    assign rom_data[1038]=8'b01101000;
    assign rom_data[1039]=8'b00111101;
    assign rom_data[1040]=8'b01101000;
    assign rom_data[1041]=8'b00111110;
    assign rom_data[1042]=8'b01101001;
    assign rom_data[1043]=8'b01000000;
    assign rom_data[1044]=8'b01101001;
    assign rom_data[1045]=8'b01000001;
    assign rom_data[1046]=8'b01101001;
    assign rom_data[1047]=8'b01000010;
    assign rom_data[1048]=8'b01101001;
    assign rom_data[1049]=8'b01000100;
    assign rom_data[1050]=8'b01101001;
    assign rom_data[1051]=8'b01000101;
    assign rom_data[1052]=8'b01101001;
    assign rom_data[1053]=8'b01000110;
    assign rom_data[1054]=8'b01101001;
    assign rom_data[1055]=8'b01000111;
    assign rom_data[1056]=8'b01101001;
    assign rom_data[1057]=8'b01001001;
    assign rom_data[1058]=8'b01101001;
    assign rom_data[1059]=8'b01001010;
    assign rom_data[1060]=8'b01101001;
    assign rom_data[1061]=8'b01001100;
    assign rom_data[1062]=8'b01101010;
    assign rom_data[1063]=8'b01001101;
    assign rom_data[1064]=8'b01101010;
    assign rom_data[1065]=8'b01001110;
    assign rom_data[1066]=8'b01101010;
    assign rom_data[1067]=8'b01010000;
    assign rom_data[1068]=8'b01101010;
    assign rom_data[1069]=8'b01010001;
    assign rom_data[1070]=8'b01101010;
    assign rom_data[1071]=8'b01010010;
    assign rom_data[1072]=8'b01101010;
    assign rom_data[1073]=8'b01010100;
    assign rom_data[1074]=8'b01101010;
    assign rom_data[1075]=8'b01010101;
    assign rom_data[1076]=8'b01101010;
    assign rom_data[1077]=8'b01010111;
    assign rom_data[1078]=8'b01101010;
    assign rom_data[1079]=8'b01011000;
    assign rom_data[1080]=8'b01101011;
    assign rom_data[1081]=8'b01011010;
    assign rom_data[1082]=8'b01101011;
    assign rom_data[1083]=8'b01011011;
    assign rom_data[1084]=8'b01101011;
    assign rom_data[1085]=8'b01011100;
    assign rom_data[1086]=8'b01101011;
    assign rom_data[1087]=8'b01011110;
    assign rom_data[1088]=8'b01101011;
    assign rom_data[1089]=8'b01011111;
    assign rom_data[1090]=8'b01101011;
    assign rom_data[1091]=8'b01100001;
    assign rom_data[1092]=8'b01101011;
    assign rom_data[1093]=8'b01100010;
    assign rom_data[1094]=8'b01101011;
    assign rom_data[1095]=8'b01100011;
    assign rom_data[1096]=8'b01101011;
    assign rom_data[1097]=8'b01100101;
    assign rom_data[1098]=8'b01101011;
    assign rom_data[1099]=8'b01100110;
    assign rom_data[1100]=8'b01101100;
    assign rom_data[1101]=8'b01100111;
    assign rom_data[1102]=8'b01101100;
    assign rom_data[1103]=8'b01101001;
    assign rom_data[1104]=8'b01101100;
    assign rom_data[1105]=8'b01101010;
    assign rom_data[1106]=8'b01101100;
    assign rom_data[1107]=8'b01101100;
    assign rom_data[1108]=8'b01101100;
    assign rom_data[1109]=8'b01101101;
    assign rom_data[1110]=8'b01101100;
    assign rom_data[1111]=8'b01101110;
    assign rom_data[1112]=8'b01101100;
    assign rom_data[1113]=8'b01110000;
    assign rom_data[1114]=8'b01101100;
    assign rom_data[1115]=8'b01110001;
    assign rom_data[1116]=8'b01101100;
    assign rom_data[1117]=8'b01110010;
    assign rom_data[1118]=8'b01101100;
    assign rom_data[1119]=8'b01110100;
    assign rom_data[1120]=8'b01101101;
    assign rom_data[1121]=8'b01110101;
    assign rom_data[1122]=8'b01101101;
    assign rom_data[1123]=8'b01110110;
    assign rom_data[1124]=8'b01101101;
    assign rom_data[1125]=8'b01110111;
    assign rom_data[1126]=8'b01101101;
    assign rom_data[1127]=8'b01111001;
    assign rom_data[1128]=8'b01101101;
    assign rom_data[1129]=8'b01111010;
    assign rom_data[1130]=8'b01101101;
    assign rom_data[1131]=8'b01111011;
    assign rom_data[1132]=8'b01101101;
    assign rom_data[1133]=8'b01111100;
    assign rom_data[1134]=8'b01101101;
    assign rom_data[1135]=8'b01111101;
    assign rom_data[1136]=8'b01101101;
    assign rom_data[1137]=8'b01111110;
    assign rom_data[1138]=8'b01101110;
    assign rom_data[1139]=8'b01111111;
    assign rom_data[1140]=8'b01101110;
    assign rom_data[1141]=8'b10000000;
    assign rom_data[1142]=8'b01101110;
    assign rom_data[1143]=8'b10000001;
    assign rom_data[1144]=8'b01101110;
    assign rom_data[1145]=8'b10000010;
    assign rom_data[1146]=8'b01101110;
    assign rom_data[1147]=8'b10000011;
    assign rom_data[1148]=8'b01101110;
    assign rom_data[1149]=8'b10000100;
    assign rom_data[1150]=8'b01101110;
    assign rom_data[1151]=8'b10000101;
    assign rom_data[1152]=8'b01101110;
    assign rom_data[1153]=8'b10000110;
    assign rom_data[1154]=8'b01101111;
    assign rom_data[1155]=8'b10000110;
    assign rom_data[1156]=8'b01101111;
    assign rom_data[1157]=8'b10000111;
    assign rom_data[1158]=8'b01101111;
    assign rom_data[1159]=8'b10001000;
    assign rom_data[1160]=8'b01101111;
    assign rom_data[1161]=8'b10001000;
    assign rom_data[1162]=8'b01101111;
    assign rom_data[1163]=8'b10001001;
    assign rom_data[1164]=8'b01101111;
    assign rom_data[1165]=8'b10001001;
    assign rom_data[1166]=8'b01101111;
    assign rom_data[1167]=8'b10001001;
    assign rom_data[1168]=8'b01110000;
    assign rom_data[1169]=8'b10001010;
    assign rom_data[1170]=8'b01110000;
    assign rom_data[1171]=8'b10001010;
    assign rom_data[1172]=8'b01110000;
    assign rom_data[1173]=8'b10001010;
    assign rom_data[1174]=8'b01110000;
    assign rom_data[1175]=8'b10001010;
    assign rom_data[1176]=8'b01110000;
    assign rom_data[1177]=8'b10001010;
    assign rom_data[1178]=8'b01110000;
    assign rom_data[1179]=8'b10001001;
    assign rom_data[1180]=8'b01110000;
    assign rom_data[1181]=8'b10001001;
    assign rom_data[1182]=8'b01110000;
    assign rom_data[1183]=8'b10001001;
    assign rom_data[1184]=8'b01110001;
    assign rom_data[1185]=8'b10001000;
    assign rom_data[1186]=8'b01110001;
    assign rom_data[1187]=8'b10001000;
    assign rom_data[1188]=8'b01110001;
    assign rom_data[1189]=8'b10000111;
    assign rom_data[1190]=8'b01110001;
    assign rom_data[1191]=8'b10000111;
    assign rom_data[1192]=8'b01110001;
    assign rom_data[1193]=8'b10000110;
    assign rom_data[1194]=8'b01110001;
    assign rom_data[1195]=8'b10000101;
    assign rom_data[1196]=8'b01110001;
    assign rom_data[1197]=8'b10000100;
    assign rom_data[1198]=8'b01110010;
    assign rom_data[1199]=8'b10000011;
    assign rom_data[1200]=8'b01110010;
    assign rom_data[1201]=8'b10000011;
    assign rom_data[1202]=8'b01110010;
    assign rom_data[1203]=8'b10000010;
    assign rom_data[1204]=8'b01110010;
    assign rom_data[1205]=8'b10000001;
    assign rom_data[1206]=8'b01110010;
    assign rom_data[1207]=8'b10000000;
    assign rom_data[1208]=8'b01110010;
    assign rom_data[1209]=8'b01111110;
    assign rom_data[1210]=8'b01110010;
    assign rom_data[1211]=8'b01111101;
    assign rom_data[1212]=8'b01110010;
    assign rom_data[1213]=8'b01111100;
    assign rom_data[1214]=8'b01110011;
    assign rom_data[1215]=8'b01111011;
    assign rom_data[1216]=8'b01110011;
    assign rom_data[1217]=8'b01111010;
    assign rom_data[1218]=8'b01110011;
    assign rom_data[1219]=8'b01111001;
    assign rom_data[1220]=8'b01110011;
    assign rom_data[1221]=8'b01110111;
    assign rom_data[1222]=8'b01110011;
    assign rom_data[1223]=8'b01110110;
    assign rom_data[1224]=8'b01110011;
    assign rom_data[1225]=8'b01110101;
    assign rom_data[1226]=8'b01110011;
    assign rom_data[1227]=8'b01110100;
    assign rom_data[1228]=8'b01110011;
    assign rom_data[1229]=8'b01110010;
    assign rom_data[1230]=8'b01110011;
    assign rom_data[1231]=8'b01110001;
    assign rom_data[1232]=8'b01110100;
    assign rom_data[1233]=8'b01110000;
    assign rom_data[1234]=8'b01110100;
    assign rom_data[1235]=8'b01101110;
    assign rom_data[1236]=8'b01110100;
    assign rom_data[1237]=8'b01101101;
    assign rom_data[1238]=8'b01110100;
    assign rom_data[1239]=8'b01101100;
    assign rom_data[1240]=8'b01110100;
    assign rom_data[1241]=8'b01101010;
    assign rom_data[1242]=8'b01110100;
    assign rom_data[1243]=8'b01101001;
    assign rom_data[1244]=8'b01110100;
    assign rom_data[1245]=8'b01100111;
    assign rom_data[1246]=8'b01110100;
    assign rom_data[1247]=8'b01100110;
    assign rom_data[1248]=8'b01110100;
    assign rom_data[1249]=8'b01100101;
    assign rom_data[1250]=8'b01110100;
    assign rom_data[1251]=8'b01100011;
    assign rom_data[1252]=8'b01110101;
    assign rom_data[1253]=8'b01100010;
    assign rom_data[1254]=8'b01110101;
    assign rom_data[1255]=8'b01100001;
    assign rom_data[1256]=8'b01110101;
    assign rom_data[1257]=8'b01011111;
    assign rom_data[1258]=8'b01110101;
    assign rom_data[1259]=8'b01011110;
    assign rom_data[1260]=8'b01110101;
    assign rom_data[1261]=8'b01011100;
    assign rom_data[1262]=8'b01110101;
    assign rom_data[1263]=8'b01011011;
    assign rom_data[1264]=8'b01110101;
    assign rom_data[1265]=8'b01011001;
    assign rom_data[1266]=8'b01110101;
    assign rom_data[1267]=8'b01011000;
    assign rom_data[1268]=8'b01110101;
    assign rom_data[1269]=8'b01010111;
    assign rom_data[1270]=8'b01110101;
    assign rom_data[1271]=8'b01010101;
    assign rom_data[1272]=8'b01110110;
    assign rom_data[1273]=8'b01010100;
    assign rom_data[1274]=8'b01110110;
    assign rom_data[1275]=8'b01010010;
    assign rom_data[1276]=8'b01110110;
    assign rom_data[1277]=8'b01010001;
    assign rom_data[1278]=8'b01110110;
    assign rom_data[1279]=8'b01010000;
    assign rom_data[1280]=8'b01110110;
    assign rom_data[1281]=8'b01001110;
    assign rom_data[1282]=8'b01110110;
    assign rom_data[1283]=8'b01001101;
    assign rom_data[1284]=8'b01110110;
    assign rom_data[1285]=8'b01001100;
    assign rom_data[1286]=8'b01110110;
    assign rom_data[1287]=8'b01001010;
    assign rom_data[1288]=8'b01110110;
    assign rom_data[1289]=8'b01001001;
    assign rom_data[1290]=8'b01110110;
    assign rom_data[1291]=8'b01001000;
    assign rom_data[1292]=8'b01110111;
    assign rom_data[1293]=8'b01000110;
    assign rom_data[1294]=8'b01110111;
    assign rom_data[1295]=8'b01000101;
    assign rom_data[1296]=8'b01110111;
    assign rom_data[1297]=8'b01000100;
    assign rom_data[1298]=8'b01110111;
    assign rom_data[1299]=8'b01000010;
    assign rom_data[1300]=8'b01110111;
    assign rom_data[1301]=8'b01000001;
    assign rom_data[1302]=8'b01110111;
    assign rom_data[1303]=8'b01000000;
    assign rom_data[1304]=8'b01110111;
    assign rom_data[1305]=8'b00111111;
    assign rom_data[1306]=8'b01110111;
    assign rom_data[1307]=8'b00111101;
    assign rom_data[1308]=8'b01110111;
    assign rom_data[1309]=8'b00111100;
    assign rom_data[1310]=8'b01111000;
    assign rom_data[1311]=8'b00111011;
    assign rom_data[1312]=8'b01111000;
    assign rom_data[1313]=8'b00111010;
    assign rom_data[1314]=8'b01111000;
    assign rom_data[1315]=8'b00111001;
    assign rom_data[1316]=8'b01111000;
    assign rom_data[1317]=8'b00111000;
    assign rom_data[1318]=8'b01111000;
    assign rom_data[1319]=8'b00110110;
    assign rom_data[1320]=8'b01111000;
    assign rom_data[1321]=8'b00110101;
    assign rom_data[1322]=8'b01111000;
    assign rom_data[1323]=8'b00110100;
    assign rom_data[1324]=8'b01111000;
    assign rom_data[1325]=8'b00110011;
    assign rom_data[1326]=8'b01111000;
    assign rom_data[1327]=8'b00110011;
    assign rom_data[1328]=8'b01111001;
    assign rom_data[1329]=8'b00110010;
    assign rom_data[1330]=8'b01111001;
    assign rom_data[1331]=8'b00110001;
    assign rom_data[1332]=8'b01111001;
    assign rom_data[1333]=8'b00110000;
    assign rom_data[1334]=8'b01111001;
    assign rom_data[1335]=8'b00101111;
    assign rom_data[1336]=8'b01111001;
    assign rom_data[1337]=8'b00101111;
    assign rom_data[1338]=8'b01111001;
    assign rom_data[1339]=8'b00101110;
    assign rom_data[1340]=8'b01111001;
    assign rom_data[1341]=8'b00101110;
    assign rom_data[1342]=8'b01111010;
    assign rom_data[1343]=8'b00101101;
    assign rom_data[1344]=8'b01111010;
    assign rom_data[1345]=8'b00101101;
    assign rom_data[1346]=8'b01111010;
    assign rom_data[1347]=8'b00101100;
    assign rom_data[1348]=8'b01111010;
    assign rom_data[1349]=8'b00101100;
    assign rom_data[1350]=8'b01111010;
    assign rom_data[1351]=8'b00101100;
    assign rom_data[1352]=8'b01111010;
    assign rom_data[1353]=8'b00101100;
    assign rom_data[1354]=8'b01111010;
    assign rom_data[1355]=8'b00101100;
    assign rom_data[1356]=8'b01111011;
    assign rom_data[1357]=8'b00101100;
    assign rom_data[1358]=8'b01111011;
    assign rom_data[1359]=8'b00101100;
    assign rom_data[1360]=8'b01111011;
    assign rom_data[1361]=8'b00101101;
    assign rom_data[1362]=8'b01111011;
    assign rom_data[1363]=8'b00101101;
    assign rom_data[1364]=8'b01111011;
    assign rom_data[1365]=8'b00101101;
    assign rom_data[1366]=8'b01111011;
    assign rom_data[1367]=8'b00101110;
    assign rom_data[1368]=8'b01111011;
    assign rom_data[1369]=8'b00101111;
    assign rom_data[1370]=8'b01111011;
    assign rom_data[1371]=8'b00101111;
    assign rom_data[1372]=8'b01111100;
    assign rom_data[1373]=8'b00110000;
    assign rom_data[1374]=8'b01111100;
    assign rom_data[1375]=8'b00110001;
    assign rom_data[1376]=8'b01111100;
    assign rom_data[1377]=8'b00110001;
    assign rom_data[1378]=8'b01111100;
    assign rom_data[1379]=8'b00110010;
    assign rom_data[1380]=8'b01111100;
    assign rom_data[1381]=8'b00110011;
    assign rom_data[1382]=8'b01111100;
    assign rom_data[1383]=8'b00110100;
    assign rom_data[1384]=8'b01111100;
    assign rom_data[1385]=8'b00110101;
    assign rom_data[1386]=8'b01111100;
    assign rom_data[1387]=8'b00110110;
    assign rom_data[1388]=8'b01111101;
    assign rom_data[1389]=8'b00110111;
    assign rom_data[1390]=8'b01111101;
    assign rom_data[1391]=8'b00111000;
    assign rom_data[1392]=8'b01111101;
    assign rom_data[1393]=8'b00111010;
    assign rom_data[1394]=8'b01111101;
    assign rom_data[1395]=8'b00111011;
    assign rom_data[1396]=8'b01111101;
    assign rom_data[1397]=8'b00111100;
    assign rom_data[1398]=8'b01111101;
    assign rom_data[1399]=8'b00111101;
    assign rom_data[1400]=8'b01111101;
    assign rom_data[1401]=8'b00111110;
    assign rom_data[1402]=8'b01111101;
    assign rom_data[1403]=8'b01000000;
    assign rom_data[1404]=8'b01111110;
    assign rom_data[1405]=8'b01000001;
    assign rom_data[1406]=8'b01111110;
    assign rom_data[1407]=8'b01000010;
    assign rom_data[1408]=8'b01111110;
    assign rom_data[1409]=8'b01000100;
    assign rom_data[1410]=8'b01111110;
    assign rom_data[1411]=8'b01000101;
    assign rom_data[1412]=8'b01111110;
    assign rom_data[1413]=8'b01000110;
    assign rom_data[1414]=8'b01111110;
    assign rom_data[1415]=8'b01000111;
    assign rom_data[1416]=8'b01111110;
    assign rom_data[1417]=8'b01001001;
    assign rom_data[1418]=8'b01111110;
    assign rom_data[1419]=8'b01001010;
    assign rom_data[1420]=8'b01111110;
    assign rom_data[1421]=8'b01001100;
    assign rom_data[1422]=8'b01111110;
    assign rom_data[1423]=8'b01001101;
    assign rom_data[1424]=8'b01111111;
    assign rom_data[1425]=8'b01001110;
    assign rom_data[1426]=8'b01111111;
    assign rom_data[1427]=8'b01010000;
    assign rom_data[1428]=8'b01111111;
    assign rom_data[1429]=8'b01010001;
    assign rom_data[1430]=8'b01111111;
    assign rom_data[1431]=8'b01010010;
    assign rom_data[1432]=8'b01111111;
    assign rom_data[1433]=8'b01010100;
    assign rom_data[1434]=8'b01111111;
    assign rom_data[1435]=8'b01010101;
    assign rom_data[1436]=8'b01111111;
    assign rom_data[1437]=8'b01010111;
    assign rom_data[1438]=8'b01111111;
    assign rom_data[1439]=8'b01011000;
    assign rom_data[1440]=8'b01111111;
    assign rom_data[1441]=8'b01011010;
    assign rom_data[1442]=8'b01111111;
    assign rom_data[1443]=8'b01011011;
    assign rom_data[1444]=8'b10000000;
    assign rom_data[1445]=8'b01011100;
    assign rom_data[1446]=8'b10000000;
    assign rom_data[1447]=8'b01011110;
    assign rom_data[1448]=8'b10000000;
    assign rom_data[1449]=8'b01011111;
    assign rom_data[1450]=8'b10000000;
    assign rom_data[1451]=8'b01100001;
    assign rom_data[1452]=8'b10000000;
    assign rom_data[1453]=8'b01100010;
    assign rom_data[1454]=8'b10000000;
    assign rom_data[1455]=8'b01100011;
    assign rom_data[1456]=8'b10000000;
    assign rom_data[1457]=8'b01100101;
    assign rom_data[1458]=8'b10000000;
    assign rom_data[1459]=8'b01100110;
    assign rom_data[1460]=8'b10000000;
    assign rom_data[1461]=8'b01100111;
    assign rom_data[1462]=8'b10000000;
    assign rom_data[1463]=8'b01101001;
    assign rom_data[1464]=8'b10000001;
    assign rom_data[1465]=8'b01101010;
    assign rom_data[1466]=8'b10000001;
    assign rom_data[1467]=8'b01101100;
    assign rom_data[1468]=8'b10000001;
    assign rom_data[1469]=8'b01101101;
    assign rom_data[1470]=8'b10000001;
    assign rom_data[1471]=8'b01101110;
    assign rom_data[1472]=8'b10000001;
    assign rom_data[1473]=8'b01110000;
    assign rom_data[1474]=8'b10000001;
    assign rom_data[1475]=8'b01110001;
    assign rom_data[1476]=8'b10000001;
    assign rom_data[1477]=8'b01110010;
    assign rom_data[1478]=8'b10000001;
    assign rom_data[1479]=8'b01110100;
    assign rom_data[1480]=8'b10000001;
    assign rom_data[1481]=8'b01110101;
    assign rom_data[1482]=8'b10000010;
    assign rom_data[1483]=8'b01110110;
    assign rom_data[1484]=8'b10000010;
    assign rom_data[1485]=8'b01110111;
    assign rom_data[1486]=8'b10000010;
    assign rom_data[1487]=8'b01111001;
    assign rom_data[1488]=8'b10000010;
    assign rom_data[1489]=8'b01111010;
    assign rom_data[1490]=8'b10000010;
    assign rom_data[1491]=8'b01111011;
    assign rom_data[1492]=8'b10000010;
    assign rom_data[1493]=8'b01111100;
    assign rom_data[1494]=8'b10000010;
    assign rom_data[1495]=8'b01111101;
    assign rom_data[1496]=8'b10000010;
    assign rom_data[1497]=8'b01111110;
    assign rom_data[1498]=8'b10000010;
    assign rom_data[1499]=8'b01111111;
    assign rom_data[1500]=8'b10000011;
    assign rom_data[1501]=8'b10000000;
    assign rom_data[1502]=8'b10000011;
    assign rom_data[1503]=8'b10000001;
    assign rom_data[1504]=8'b10000011;
    assign rom_data[1505]=8'b10000010;
    assign rom_data[1506]=8'b10000011;
    assign rom_data[1507]=8'b10000011;
    assign rom_data[1508]=8'b10000011;
    assign rom_data[1509]=8'b10000100;
    assign rom_data[1510]=8'b10000011;
    assign rom_data[1511]=8'b10000101;
    assign rom_data[1512]=8'b10000011;
    assign rom_data[1513]=8'b10000110;
    assign rom_data[1514]=8'b10000011;
    assign rom_data[1515]=8'b10000110;
    assign rom_data[1516]=8'b10000100;
    assign rom_data[1517]=8'b10000111;
    assign rom_data[1518]=8'b10000100;
    assign rom_data[1519]=8'b10001000;
    assign rom_data[1520]=8'b10000100;
    assign rom_data[1521]=8'b10001000;
    assign rom_data[1522]=8'b10000100;
    assign rom_data[1523]=8'b10001001;
    assign rom_data[1524]=8'b10000100;
    assign rom_data[1525]=8'b10001001;
    assign rom_data[1526]=8'b10000100;
    assign rom_data[1527]=8'b10001001;
    assign rom_data[1528]=8'b10000100;
    assign rom_data[1529]=8'b10001010;
    assign rom_data[1530]=8'b10000101;
    assign rom_data[1531]=8'b10001010;
    assign rom_data[1532]=8'b10000101;
    assign rom_data[1533]=8'b10001010;
    assign rom_data[1534]=8'b10000101;
    assign rom_data[1535]=8'b10001010;
    assign rom_data[1536]=8'b10000101;
    assign rom_data[1537]=8'b10001010;
    assign rom_data[1538]=8'b10000101;
    assign rom_data[1539]=8'b10001001;
    assign rom_data[1540]=8'b10000101;
    assign rom_data[1541]=8'b10001001;
    assign rom_data[1542]=8'b10000101;
    assign rom_data[1543]=8'b10001001;
    assign rom_data[1544]=8'b10000101;
    assign rom_data[1545]=8'b10001000;
    assign rom_data[1546]=8'b10000110;
    assign rom_data[1547]=8'b10001000;
    assign rom_data[1548]=8'b10000110;
    assign rom_data[1549]=8'b10000111;
    assign rom_data[1550]=8'b10000110;
    assign rom_data[1551]=8'b10000111;
    assign rom_data[1552]=8'b10000110;
    assign rom_data[1553]=8'b10000110;
    assign rom_data[1554]=8'b10000110;
    assign rom_data[1555]=8'b10000101;
    assign rom_data[1556]=8'b10000110;
    assign rom_data[1557]=8'b10000100;
    assign rom_data[1558]=8'b10000110;
    assign rom_data[1559]=8'b10000011;
    assign rom_data[1560]=8'b10000111;
    assign rom_data[1561]=8'b10000011;
    assign rom_data[1562]=8'b10000111;
    assign rom_data[1563]=8'b10000010;
    assign rom_data[1564]=8'b10000111;
    assign rom_data[1565]=8'b10000001;
    assign rom_data[1566]=8'b10000111;
    assign rom_data[1567]=8'b10000000;
    assign rom_data[1568]=8'b10000111;
    assign rom_data[1569]=8'b01111110;
    assign rom_data[1570]=8'b10000111;
    assign rom_data[1571]=8'b01111101;
    assign rom_data[1572]=8'b10000111;
    assign rom_data[1573]=8'b01111100;
    assign rom_data[1574]=8'b10000111;
    assign rom_data[1575]=8'b01111011;
    assign rom_data[1576]=8'b10000111;
    assign rom_data[1577]=8'b01111010;
    assign rom_data[1578]=8'b10001000;
    assign rom_data[1579]=8'b01111001;
    assign rom_data[1580]=8'b10001000;
    assign rom_data[1581]=8'b01110111;
    assign rom_data[1582]=8'b10001000;
    assign rom_data[1583]=8'b01110110;
    assign rom_data[1584]=8'b10001000;
    assign rom_data[1585]=8'b01110101;
    assign rom_data[1586]=8'b10001000;
    assign rom_data[1587]=8'b01110100;
    assign rom_data[1588]=8'b10001000;
    assign rom_data[1589]=8'b01110010;
    assign rom_data[1590]=8'b10001000;
    assign rom_data[1591]=8'b01110001;
    assign rom_data[1592]=8'b10001000;
    assign rom_data[1593]=8'b01110000;
    assign rom_data[1594]=8'b10001000;
    assign rom_data[1595]=8'b01101110;
    assign rom_data[1596]=8'b10001001;
    assign rom_data[1597]=8'b01101101;
    assign rom_data[1598]=8'b10001001;
    assign rom_data[1599]=8'b01101100;
    assign rom_data[1600]=8'b10001001;
    assign rom_data[1601]=8'b01101010;
    assign rom_data[1602]=8'b10001001;
    assign rom_data[1603]=8'b01101001;
    assign rom_data[1604]=8'b10001001;
    assign rom_data[1605]=8'b01100111;
    assign rom_data[1606]=8'b10001001;
    assign rom_data[1607]=8'b01100110;
    assign rom_data[1608]=8'b10001001;
    assign rom_data[1609]=8'b01100101;
    assign rom_data[1610]=8'b10001001;
    assign rom_data[1611]=8'b01100011;
    assign rom_data[1612]=8'b10001001;
    assign rom_data[1613]=8'b01100010;
    assign rom_data[1614]=8'b10001001;
    assign rom_data[1615]=8'b01100001;
    assign rom_data[1616]=8'b10001010;
    assign rom_data[1617]=8'b01011111;
    assign rom_data[1618]=8'b10001010;
    assign rom_data[1619]=8'b01011110;
    assign rom_data[1620]=8'b10001010;
    assign rom_data[1621]=8'b01011100;
    assign rom_data[1622]=8'b10001010;
    assign rom_data[1623]=8'b01011011;
    assign rom_data[1624]=8'b10001010;
    assign rom_data[1625]=8'b01011001;
    assign rom_data[1626]=8'b10001010;
    assign rom_data[1627]=8'b01011000;
    assign rom_data[1628]=8'b10001001;
    assign rom_data[1629]=8'b01010111;
    assign rom_data[1630]=8'b10001001;
    assign rom_data[1631]=8'b01010101;
    assign rom_data[1632]=8'b10001001;
    assign rom_data[1633]=8'b01010100;
    assign rom_data[1634]=8'b10001001;
    assign rom_data[1635]=8'b01010010;
    assign rom_data[1636]=8'b10001001;
    assign rom_data[1637]=8'b01010001;
    assign rom_data[1638]=8'b10001001;
    assign rom_data[1639]=8'b01010000;
    assign rom_data[1640]=8'b10001001;
    assign rom_data[1641]=8'b01001110;
    assign rom_data[1642]=8'b10001001;
    assign rom_data[1643]=8'b01001101;
    assign rom_data[1644]=8'b10001001;
    assign rom_data[1645]=8'b01001100;
    assign rom_data[1646]=8'b10001001;
    assign rom_data[1647]=8'b01001010;
    assign rom_data[1648]=8'b10001000;
    assign rom_data[1649]=8'b01001001;
    assign rom_data[1650]=8'b10001000;
    assign rom_data[1651]=8'b01001000;
    assign rom_data[1652]=8'b10001000;
    assign rom_data[1653]=8'b01000110;
    assign rom_data[1654]=8'b10001000;
    assign rom_data[1655]=8'b01000101;
    assign rom_data[1656]=8'b10001000;
    assign rom_data[1657]=8'b01000100;
    assign rom_data[1658]=8'b10001000;
    assign rom_data[1659]=8'b01000010;
    assign rom_data[1660]=8'b10001000;
    assign rom_data[1661]=8'b01000001;
    assign rom_data[1662]=8'b10001000;
    assign rom_data[1663]=8'b01000000;
    assign rom_data[1664]=8'b10001000;
    assign rom_data[1665]=8'b00111111;
    assign rom_data[1666]=8'b10000111;
    assign rom_data[1667]=8'b00111101;
    assign rom_data[1668]=8'b10000111;
    assign rom_data[1669]=8'b00111100;
    assign rom_data[1670]=8'b10000111;
    assign rom_data[1671]=8'b00111011;
    assign rom_data[1672]=8'b10000111;
    assign rom_data[1673]=8'b00111010;
    assign rom_data[1674]=8'b10000111;
    assign rom_data[1675]=8'b00111001;
    assign rom_data[1676]=8'b10000111;
    assign rom_data[1677]=8'b00111000;
    assign rom_data[1678]=8'b10000111;
    assign rom_data[1679]=8'b00110110;
    assign rom_data[1680]=8'b10000111;
    assign rom_data[1681]=8'b00110101;
    assign rom_data[1682]=8'b10000111;
    assign rom_data[1683]=8'b00110100;
    assign rom_data[1684]=8'b10000110;
    assign rom_data[1685]=8'b00110011;
    assign rom_data[1686]=8'b10000110;
    assign rom_data[1687]=8'b00110011;
    assign rom_data[1688]=8'b10000110;
    assign rom_data[1689]=8'b00110010;
    assign rom_data[1690]=8'b10000110;
    assign rom_data[1691]=8'b00110001;
    assign rom_data[1692]=8'b10000110;
    assign rom_data[1693]=8'b00110000;
    assign rom_data[1694]=8'b10000110;
    assign rom_data[1695]=8'b00101111;
    assign rom_data[1696]=8'b10000110;
    assign rom_data[1697]=8'b00101111;
    assign rom_data[1698]=8'b10000101;
    assign rom_data[1699]=8'b00101110;
    assign rom_data[1700]=8'b10000101;
    assign rom_data[1701]=8'b00101110;
    assign rom_data[1702]=8'b10000101;
    assign rom_data[1703]=8'b00101101;
    assign rom_data[1704]=8'b10000101;
    assign rom_data[1705]=8'b00101101;
    assign rom_data[1706]=8'b10000101;
    assign rom_data[1707]=8'b00101100;
    assign rom_data[1708]=8'b10000101;
    assign rom_data[1709]=8'b00101100;
    assign rom_data[1710]=8'b10000101;
    assign rom_data[1711]=8'b00101100;
    assign rom_data[1712]=8'b10000101;
    assign rom_data[1713]=8'b00101100;
    assign rom_data[1714]=8'b10000100;
    assign rom_data[1715]=8'b00101100;
    assign rom_data[1716]=8'b10000100;
    assign rom_data[1717]=8'b00101100;
    assign rom_data[1718]=8'b10000100;
    assign rom_data[1719]=8'b00101100;
    assign rom_data[1720]=8'b10000100;
    assign rom_data[1721]=8'b00101101;
    assign rom_data[1722]=8'b10000100;
    assign rom_data[1723]=8'b00101101;
    assign rom_data[1724]=8'b10000100;
    assign rom_data[1725]=8'b00101101;
    assign rom_data[1726]=8'b10000100;
    assign rom_data[1727]=8'b00101110;
    assign rom_data[1728]=8'b10000011;
    assign rom_data[1729]=8'b00101111;
    assign rom_data[1730]=8'b10000011;
    assign rom_data[1731]=8'b00101111;
    assign rom_data[1732]=8'b10000011;
    assign rom_data[1733]=8'b00110000;
    assign rom_data[1734]=8'b10000011;
    assign rom_data[1735]=8'b00110001;
    assign rom_data[1736]=8'b10000011;
    assign rom_data[1737]=8'b00110001;
    assign rom_data[1738]=8'b10000011;
    assign rom_data[1739]=8'b00110010;
    assign rom_data[1740]=8'b10000011;
    assign rom_data[1741]=8'b00110011;
    assign rom_data[1742]=8'b10000011;
    assign rom_data[1743]=8'b00110100;
    assign rom_data[1744]=8'b10000010;
    assign rom_data[1745]=8'b00110101;
    assign rom_data[1746]=8'b10000010;
    assign rom_data[1747]=8'b00110110;
    assign rom_data[1748]=8'b10000010;
    assign rom_data[1749]=8'b00110111;
    assign rom_data[1750]=8'b10000010;
    assign rom_data[1751]=8'b00111000;
    assign rom_data[1752]=8'b10000010;
    assign rom_data[1753]=8'b00111010;
    assign rom_data[1754]=8'b10000010;
    assign rom_data[1755]=8'b00111011;
    assign rom_data[1756]=8'b10000010;
    assign rom_data[1757]=8'b00111100;
    assign rom_data[1758]=8'b10000010;
    assign rom_data[1759]=8'b00111101;
    assign rom_data[1760]=8'b10000010;
    assign rom_data[1761]=8'b00111110;
    assign rom_data[1762]=8'b10000001;
    assign rom_data[1763]=8'b01000000;
    assign rom_data[1764]=8'b10000001;
    assign rom_data[1765]=8'b01000001;
    assign rom_data[1766]=8'b10000001;
    assign rom_data[1767]=8'b01000010;
    assign rom_data[1768]=8'b10000001;
    assign rom_data[1769]=8'b01000100;
    assign rom_data[1770]=8'b10000001;
    assign rom_data[1771]=8'b01000101;
    assign rom_data[1772]=8'b10000001;
    assign rom_data[1773]=8'b01000110;
    assign rom_data[1774]=8'b10000001;
    assign rom_data[1775]=8'b01000111;
    assign rom_data[1776]=8'b10000001;
    assign rom_data[1777]=8'b01001001;
    assign rom_data[1778]=8'b10000001;
    assign rom_data[1779]=8'b01001010;
    assign rom_data[1780]=8'b10000000;
    assign rom_data[1781]=8'b01001100;
    assign rom_data[1782]=8'b10000000;
    assign rom_data[1783]=8'b01001101;
    assign rom_data[1784]=8'b10000000;
    assign rom_data[1785]=8'b01001110;
    assign rom_data[1786]=8'b10000000;
    assign rom_data[1787]=8'b01010000;
    assign rom_data[1788]=8'b10000000;
    assign rom_data[1789]=8'b01010001;
    assign rom_data[1790]=8'b10000000;
    assign rom_data[1791]=8'b01010010;
    assign rom_data[1792]=8'b10000000;
    assign rom_data[1793]=8'b01010100;
    assign rom_data[1794]=8'b10000000;
    assign rom_data[1795]=8'b01010101;
    assign rom_data[1796]=8'b10000000;
    assign rom_data[1797]=8'b01010111;
    assign rom_data[1798]=8'b10000000;
    assign rom_data[1799]=8'b01011000;
    assign rom_data[1800]=8'b01111111;
    assign rom_data[1801]=8'b01011010;
    assign rom_data[1802]=8'b01111111;
    assign rom_data[1803]=8'b01011011;
    assign rom_data[1804]=8'b01111111;
    assign rom_data[1805]=8'b01011100;
    assign rom_data[1806]=8'b01111111;
    assign rom_data[1807]=8'b01011110;
    assign rom_data[1808]=8'b01111111;
    assign rom_data[1809]=8'b01011111;
    assign rom_data[1810]=8'b01111111;
    assign rom_data[1811]=8'b01100001;
    assign rom_data[1812]=8'b01111111;
    assign rom_data[1813]=8'b01100010;
    assign rom_data[1814]=8'b01111111;
    assign rom_data[1815]=8'b01100011;
    assign rom_data[1816]=8'b01111111;
    assign rom_data[1817]=8'b01100101;
    assign rom_data[1818]=8'b01111111;
    assign rom_data[1819]=8'b01100110;
    assign rom_data[1820]=8'b01111110;
    assign rom_data[1821]=8'b01100111;
    assign rom_data[1822]=8'b01111110;
    assign rom_data[1823]=8'b01101001;
    assign rom_data[1824]=8'b01111110;
    assign rom_data[1825]=8'b01101010;
    assign rom_data[1826]=8'b01111110;
    assign rom_data[1827]=8'b01101100;
    assign rom_data[1828]=8'b01111110;
    assign rom_data[1829]=8'b01101101;
    assign rom_data[1830]=8'b01111110;
    assign rom_data[1831]=8'b01101110;
    assign rom_data[1832]=8'b01111110;
    assign rom_data[1833]=8'b01110000;
    assign rom_data[1834]=8'b01111110;
    assign rom_data[1835]=8'b01110001;
    assign rom_data[1836]=8'b01111110;
    assign rom_data[1837]=8'b01110010;
    assign rom_data[1838]=8'b01111110;
    assign rom_data[1839]=8'b01110100;
    assign rom_data[1840]=8'b01111101;
    assign rom_data[1841]=8'b01110101;
    assign rom_data[1842]=8'b01111101;
    assign rom_data[1843]=8'b01110110;
    assign rom_data[1844]=8'b01111101;
    assign rom_data[1845]=8'b01110111;
    assign rom_data[1846]=8'b01111101;
    assign rom_data[1847]=8'b01111001;
    assign rom_data[1848]=8'b01111101;
    assign rom_data[1849]=8'b01111010;
    assign rom_data[1850]=8'b01111101;
    assign rom_data[1851]=8'b01111011;
    assign rom_data[1852]=8'b01111101;
    assign rom_data[1853]=8'b01111100;
    assign rom_data[1854]=8'b01111101;
    assign rom_data[1855]=8'b01111101;
    assign rom_data[1856]=8'b01111100;
    assign rom_data[1857]=8'b01111110;
    assign rom_data[1858]=8'b01111100;
    assign rom_data[1859]=8'b01111111;
    assign rom_data[1860]=8'b01111100;
    assign rom_data[1861]=8'b10000000;
    assign rom_data[1862]=8'b01111100;
    assign rom_data[1863]=8'b10000001;
    assign rom_data[1864]=8'b01111100;
    assign rom_data[1865]=8'b10000010;
    assign rom_data[1866]=8'b01111100;
    assign rom_data[1867]=8'b10000011;
    assign rom_data[1868]=8'b01111100;
    assign rom_data[1869]=8'b10000100;
    assign rom_data[1870]=8'b01111100;
    assign rom_data[1871]=8'b10000101;
    assign rom_data[1872]=8'b01111011;
    assign rom_data[1873]=8'b10000110;
    assign rom_data[1874]=8'b01111011;
    assign rom_data[1875]=8'b10000110;
    assign rom_data[1876]=8'b01111011;
    assign rom_data[1877]=8'b10000111;
    assign rom_data[1878]=8'b01111011;
    assign rom_data[1879]=8'b10001000;
    assign rom_data[1880]=8'b01111011;
    assign rom_data[1881]=8'b10001000;
    assign rom_data[1882]=8'b01111011;
    assign rom_data[1883]=8'b10001001;
    assign rom_data[1884]=8'b01111011;
    assign rom_data[1885]=8'b10001001;
    assign rom_data[1886]=8'b01111011;
    assign rom_data[1887]=8'b10001001;
    assign rom_data[1888]=8'b01111010;
    assign rom_data[1889]=8'b10001010;
    assign rom_data[1890]=8'b01111010;
    assign rom_data[1891]=8'b10001010;
    assign rom_data[1892]=8'b01111010;
    assign rom_data[1893]=8'b10001010;
    assign rom_data[1894]=8'b01111010;
    assign rom_data[1895]=8'b10001010;
    assign rom_data[1896]=8'b01111010;
    assign rom_data[1897]=8'b10001010;
    assign rom_data[1898]=8'b01111010;
    assign rom_data[1899]=8'b10001001;
    assign rom_data[1900]=8'b01111010;
    assign rom_data[1901]=8'b10001001;
    assign rom_data[1902]=8'b01111001;
    assign rom_data[1903]=8'b10001001;
    assign rom_data[1904]=8'b01111001;
    assign rom_data[1905]=8'b10001000;
    assign rom_data[1906]=8'b01111001;
    assign rom_data[1907]=8'b10001000;
    assign rom_data[1908]=8'b01111001;
    assign rom_data[1909]=8'b10000111;
    assign rom_data[1910]=8'b01111001;
    assign rom_data[1911]=8'b10000111;
    assign rom_data[1912]=8'b01111001;
    assign rom_data[1913]=8'b10000110;
    assign rom_data[1914]=8'b01111001;
    assign rom_data[1915]=8'b10000101;
    assign rom_data[1916]=8'b01111000;
    assign rom_data[1917]=8'b10000100;
    assign rom_data[1918]=8'b01111000;
    assign rom_data[1919]=8'b10000011;
    assign rom_data[1920]=8'b01111000;
    assign rom_data[1921]=8'b10000011;
    assign rom_data[1922]=8'b01111000;
    assign rom_data[1923]=8'b10000010;
    assign rom_data[1924]=8'b01111000;
    assign rom_data[1925]=8'b10000001;
    assign rom_data[1926]=8'b01111000;
    assign rom_data[1927]=8'b10000000;
    assign rom_data[1928]=8'b01111000;
    assign rom_data[1929]=8'b01111110;
    assign rom_data[1930]=8'b01111000;
    assign rom_data[1931]=8'b01111101;
    assign rom_data[1932]=8'b01111000;
    assign rom_data[1933]=8'b01111100;
    assign rom_data[1934]=8'b01110111;
    assign rom_data[1935]=8'b01111011;
    assign rom_data[1936]=8'b01110111;
    assign rom_data[1937]=8'b01111010;
    assign rom_data[1938]=8'b01110111;
    assign rom_data[1939]=8'b01111001;
    assign rom_data[1940]=8'b01110111;
    assign rom_data[1941]=8'b01110111;
    assign rom_data[1942]=8'b01110111;
    assign rom_data[1943]=8'b01110110;
    assign rom_data[1944]=8'b01110111;
    assign rom_data[1945]=8'b01110101;
    assign rom_data[1946]=8'b01110111;
    assign rom_data[1947]=8'b01110100;
    assign rom_data[1948]=8'b01110111;
    assign rom_data[1949]=8'b01110010;
    assign rom_data[1950]=8'b01110111;
    assign rom_data[1951]=8'b01110001;
    assign rom_data[1952]=8'b01110110;
    assign rom_data[1953]=8'b01110000;
    assign rom_data[1954]=8'b01110110;
    assign rom_data[1955]=8'b01101110;
    assign rom_data[1956]=8'b01110110;
    assign rom_data[1957]=8'b01101101;
    assign rom_data[1958]=8'b01110110;
    assign rom_data[1959]=8'b01101100;
    assign rom_data[1960]=8'b01110110;
    assign rom_data[1961]=8'b01101010;
    assign rom_data[1962]=8'b01110110;
    assign rom_data[1963]=8'b01101001;
    assign rom_data[1964]=8'b01110110;
    assign rom_data[1965]=8'b01100111;
    assign rom_data[1966]=8'b01110110;
    assign rom_data[1967]=8'b01100110;
    assign rom_data[1968]=8'b01110110;
    assign rom_data[1969]=8'b01100101;
    assign rom_data[1970]=8'b01110110;
    assign rom_data[1971]=8'b01100011;
    assign rom_data[1972]=8'b01110101;
    assign rom_data[1973]=8'b01100010;
    assign rom_data[1974]=8'b01110101;
    assign rom_data[1975]=8'b01100001;
    assign rom_data[1976]=8'b01110101;
    assign rom_data[1977]=8'b01011111;
    assign rom_data[1978]=8'b01110101;
    assign rom_data[1979]=8'b01011110;
    assign rom_data[1980]=8'b01110101;
    assign rom_data[1981]=8'b01011100;
    assign rom_data[1982]=8'b01110101;
    assign rom_data[1983]=8'b01011011;
    assign rom_data[1984]=8'b01110101;
    assign rom_data[1985]=8'b01011001;
    assign rom_data[1986]=8'b01110101;
    assign rom_data[1987]=8'b01011000;
    assign rom_data[1988]=8'b01110101;
    assign rom_data[1989]=8'b01010111;
    assign rom_data[1990]=8'b01110101;
    assign rom_data[1991]=8'b01010101;
    assign rom_data[1992]=8'b01110100;
    assign rom_data[1993]=8'b01010100;
    assign rom_data[1994]=8'b01110100;
    assign rom_data[1995]=8'b01010010;
    assign rom_data[1996]=8'b01110100;
    assign rom_data[1997]=8'b01010001;
    assign rom_data[1998]=8'b01110100;
    assign rom_data[1999]=8'b01010000;
    assign rom_data[2000]=8'b01110100;
    assign rom_data[2001]=8'b01001110;
    assign rom_data[2002]=8'b01110100;
    assign rom_data[2003]=8'b01001101;
    assign rom_data[2004]=8'b01110100;
    assign rom_data[2005]=8'b01001100;
    assign rom_data[2006]=8'b01110100;
    assign rom_data[2007]=8'b01001010;
    assign rom_data[2008]=8'b01110100;
    assign rom_data[2009]=8'b01001001;
    assign rom_data[2010]=8'b01110100;
    assign rom_data[2011]=8'b01001000;
    assign rom_data[2012]=8'b01110011;
    assign rom_data[2013]=8'b01000110;
    assign rom_data[2014]=8'b01110011;
    assign rom_data[2015]=8'b01000101;
    assign rom_data[2016]=8'b01110011;
    assign rom_data[2017]=8'b01000100;
    assign rom_data[2018]=8'b01110011;
    assign rom_data[2019]=8'b01000010;
    assign rom_data[2020]=8'b01110011;
    assign rom_data[2021]=8'b01000001;
    assign rom_data[2022]=8'b01110011;
    assign rom_data[2023]=8'b01000000;
    assign rom_data[2024]=8'b01110011;
    assign rom_data[2025]=8'b00111111;
    assign rom_data[2026]=8'b01110011;
    assign rom_data[2027]=8'b00111101;
    assign rom_data[2028]=8'b01110011;
    assign rom_data[2029]=8'b00111100;
    assign rom_data[2030]=8'b01110010;
    assign rom_data[2031]=8'b00111011;
    assign rom_data[2032]=8'b01110010;
    assign rom_data[2033]=8'b00111010;
    assign rom_data[2034]=8'b01110010;
    assign rom_data[2035]=8'b00111001;
    assign rom_data[2036]=8'b01110010;
    assign rom_data[2037]=8'b00111000;
    assign rom_data[2038]=8'b01110010;
    assign rom_data[2039]=8'b00110110;
    assign rom_data[2040]=8'b01110010;
    assign rom_data[2041]=8'b00110101;
    assign rom_data[2042]=8'b01110010;
    assign rom_data[2043]=8'b00110100;
    assign rom_data[2044]=8'b01110010;
    assign rom_data[2045]=8'b00110011;
    assign rom_data[2046]=8'b01110001;
    assign rom_data[2047]=8'b00110011;
    assign rom_data[2048]=8'b01110001;
    assign rom_data[2049]=8'b00110010;
    assign rom_data[2050]=8'b01110001;
    assign rom_data[2051]=8'b00110001;
    assign rom_data[2052]=8'b01110001;
    assign rom_data[2053]=8'b00110000;
    assign rom_data[2054]=8'b01110001;
    assign rom_data[2055]=8'b00101111;
    assign rom_data[2056]=8'b01110001;
    assign rom_data[2057]=8'b00101111;
    assign rom_data[2058]=8'b01110001;
    assign rom_data[2059]=8'b00101110;
    assign rom_data[2060]=8'b01110000;
    assign rom_data[2061]=8'b00101110;
    assign rom_data[2062]=8'b01110000;
    assign rom_data[2063]=8'b00101101;
    assign rom_data[2064]=8'b01110000;
    assign rom_data[2065]=8'b00101101;
    assign rom_data[2066]=8'b01110000;
    assign rom_data[2067]=8'b00101100;
    assign rom_data[2068]=8'b01110000;
    assign rom_data[2069]=8'b00101100;
    assign rom_data[2070]=8'b01110000;
    assign rom_data[2071]=8'b00101100;
    assign rom_data[2072]=8'b01110000;
    assign rom_data[2073]=8'b00101100;
    assign rom_data[2074]=8'b01110000;
    assign rom_data[2075]=8'b00101100;
    assign rom_data[2076]=8'b01101111;
    assign rom_data[2077]=8'b00101100;
    assign rom_data[2078]=8'b01101111;
    assign rom_data[2079]=8'b00101100;
    assign rom_data[2080]=8'b01101111;
    assign rom_data[2081]=8'b00101101;
    assign rom_data[2082]=8'b01101111;
    assign rom_data[2083]=8'b00101101;
    assign rom_data[2084]=8'b01101111;
    assign rom_data[2085]=8'b00101101;
    assign rom_data[2086]=8'b01101111;
    assign rom_data[2087]=8'b00101110;
    assign rom_data[2088]=8'b01101111;
    assign rom_data[2089]=8'b00101111;
    assign rom_data[2090]=8'b01101110;
    assign rom_data[2091]=8'b00101111;
    assign rom_data[2092]=8'b01101110;
    assign rom_data[2093]=8'b00110000;
    assign rom_data[2094]=8'b01101110;
    assign rom_data[2095]=8'b00110001;
    assign rom_data[2096]=8'b01101110;
    assign rom_data[2097]=8'b00110001;
    assign rom_data[2098]=8'b01101110;
    assign rom_data[2099]=8'b00110010;
    assign rom_data[2100]=8'b01101110;
    assign rom_data[2101]=8'b00110011;
    assign rom_data[2102]=8'b01101110;
    assign rom_data[2103]=8'b00110100;
    assign rom_data[2104]=8'b01101110;
    assign rom_data[2105]=8'b00110101;
    assign rom_data[2106]=8'b01101101;
    assign rom_data[2107]=8'b00110110;
    assign rom_data[2108]=8'b01101101;
    assign rom_data[2109]=8'b00110111;
    assign rom_data[2110]=8'b01101101;
    assign rom_data[2111]=8'b00111000;
    assign rom_data[2112]=8'b01101101;
    assign rom_data[2113]=8'b00111010;
    assign rom_data[2114]=8'b01101101;
    assign rom_data[2115]=8'b00111011;
    assign rom_data[2116]=8'b01101101;
    assign rom_data[2117]=8'b00111100;
    assign rom_data[2118]=8'b01101101;
    assign rom_data[2119]=8'b00111101;
    assign rom_data[2120]=8'b01101101;
    assign rom_data[2121]=8'b00111110;
    assign rom_data[2122]=8'b01101101;
    assign rom_data[2123]=8'b01000000;
    assign rom_data[2124]=8'b01101100;
    assign rom_data[2125]=8'b01000001;
    assign rom_data[2126]=8'b01101100;
    assign rom_data[2127]=8'b01000010;
    assign rom_data[2128]=8'b01101100;
    assign rom_data[2129]=8'b01000100;
    assign rom_data[2130]=8'b01101100;
    assign rom_data[2131]=8'b01000101;
    assign rom_data[2132]=8'b01101100;
    assign rom_data[2133]=8'b01000110;
    assign rom_data[2134]=8'b01101100;
    assign rom_data[2135]=8'b01000111;
    assign rom_data[2136]=8'b01101100;
    assign rom_data[2137]=8'b01001001;
    assign rom_data[2138]=8'b01101100;
    assign rom_data[2139]=8'b01001010;
    assign rom_data[2140]=8'b01101100;
    assign rom_data[2141]=8'b01001100;
    assign rom_data[2142]=8'b01101100;
    assign rom_data[2143]=8'b01001101;
    assign rom_data[2144]=8'b01101011;
    assign rom_data[2145]=8'b01001110;
    assign rom_data[2146]=8'b01101011;
    assign rom_data[2147]=8'b01010000;
    assign rom_data[2148]=8'b01101011;
    assign rom_data[2149]=8'b01010001;
    assign rom_data[2150]=8'b01101011;
    assign rom_data[2151]=8'b01010010;
    assign rom_data[2152]=8'b01101011;
    assign rom_data[2153]=8'b01010100;
    assign rom_data[2154]=8'b01101011;
    assign rom_data[2155]=8'b01010101;
    assign rom_data[2156]=8'b01101011;
    assign rom_data[2157]=8'b01010111;
    assign rom_data[2158]=8'b01101011;
    assign rom_data[2159]=8'b01011000;
    assign rom_data[2160]=8'b01101011;
    assign rom_data[2161]=8'b01011010;
    assign rom_data[2162]=8'b01101011;
    assign rom_data[2163]=8'b01011011;
    assign rom_data[2164]=8'b01101010;
    assign rom_data[2165]=8'b01011100;
    assign rom_data[2166]=8'b01101010;
    assign rom_data[2167]=8'b01011110;
    assign rom_data[2168]=8'b01101010;
    assign rom_data[2169]=8'b01011111;
    assign rom_data[2170]=8'b01101010;
    assign rom_data[2171]=8'b01100001;
    assign rom_data[2172]=8'b01101010;
    assign rom_data[2173]=8'b01100010;
    assign rom_data[2174]=8'b01101010;
    assign rom_data[2175]=8'b01100011;
    assign rom_data[2176]=8'b01101010;
    assign rom_data[2177]=8'b01100101;
    assign rom_data[2178]=8'b01101010;
    assign rom_data[2179]=8'b01100110;
    assign rom_data[2180]=8'b01101010;
    assign rom_data[2181]=8'b01100111;
    assign rom_data[2182]=8'b01101001;
    assign rom_data[2183]=8'b01101001;
    assign rom_data[2184]=8'b01101001;
    assign rom_data[2185]=8'b01101010;
    assign rom_data[2186]=8'b01101001;
    assign rom_data[2187]=8'b01101100;
    assign rom_data[2188]=8'b01101001;
    assign rom_data[2189]=8'b01101101;
    assign rom_data[2190]=8'b01101001;
    assign rom_data[2191]=8'b01101110;
    assign rom_data[2192]=8'b01101001;
    assign rom_data[2193]=8'b01110000;
    assign rom_data[2194]=8'b01101001;
    assign rom_data[2195]=8'b01110001;
    assign rom_data[2196]=8'b01101001;
    assign rom_data[2197]=8'b01110010;
    assign rom_data[2198]=8'b01101001;
    assign rom_data[2199]=8'b01110100;
    assign rom_data[2200]=8'b01101001;
    assign rom_data[2201]=8'b01110101;
    assign rom_data[2202]=8'b01101000;
    assign rom_data[2203]=8'b01110110;
    assign rom_data[2204]=8'b01101000;
    assign rom_data[2205]=8'b01110111;
    assign rom_data[2206]=8'b01101000;
    assign rom_data[2207]=8'b01111001;
    assign rom_data[2208]=8'b01101000;
    assign rom_data[2209]=8'b01111010;
    assign rom_data[2210]=8'b01101000;
    assign rom_data[2211]=8'b01111011;
    assign rom_data[2212]=8'b01101000;
    assign rom_data[2213]=8'b01111100;
    assign rom_data[2214]=8'b01101000;
    assign rom_data[2215]=8'b01111101;
    assign rom_data[2216]=8'b01101000;
    assign rom_data[2217]=8'b01111110;
    assign rom_data[2218]=8'b01101000;
    assign rom_data[2219]=8'b01111111;
    assign rom_data[2220]=8'b01100111;
    assign rom_data[2221]=8'b10000000;
    assign rom_data[2222]=8'b01100111;
    assign rom_data[2223]=8'b10000001;
    assign rom_data[2224]=8'b01100111;
    assign rom_data[2225]=8'b10000010;
    assign rom_data[2226]=8'b01100111;
    assign rom_data[2227]=8'b10000011;
    assign rom_data[2228]=8'b01100111;
    assign rom_data[2229]=8'b10000100;
    assign rom_data[2230]=8'b01100111;
    assign rom_data[2231]=8'b10000101;
    assign rom_data[2232]=8'b01100111;
    assign rom_data[2233]=8'b10000110;
    assign rom_data[2234]=8'b01100110;
    assign rom_data[2235]=8'b10000110;
    assign rom_data[2236]=8'b01100110;
    assign rom_data[2237]=8'b10000111;
    assign rom_data[2238]=8'b01100110;
    assign rom_data[2239]=8'b10001000;
    assign rom_data[2240]=8'b01100110;
    assign rom_data[2241]=8'b10001000;
    assign rom_data[2242]=8'b01100110;
    assign rom_data[2243]=8'b10001001;
    assign rom_data[2244]=8'b01100110;
    assign rom_data[2245]=8'b10001001;
    assign rom_data[2246]=8'b01100110;
    assign rom_data[2247]=8'b10001001;
    assign rom_data[2248]=8'b01100110;
    assign rom_data[2249]=8'b10001010;
    assign rom_data[2250]=8'b01100101;
    assign rom_data[2251]=8'b10001010;
    assign rom_data[2252]=8'b01100101;
    assign rom_data[2253]=8'b10001010;
    assign rom_data[2254]=8'b01100101;
    assign rom_data[2255]=8'b10001010;
    assign rom_data[2256]=8'b01100101;
    assign rom_data[2257]=8'b10001010;
    assign rom_data[2258]=8'b01100101;
    assign rom_data[2259]=8'b10001001;
    assign rom_data[2260]=8'b01100101;
    assign rom_data[2261]=8'b10001001;
    assign rom_data[2262]=8'b01100101;
    assign rom_data[2263]=8'b10001001;
    assign rom_data[2264]=8'b01100100;
    assign rom_data[2265]=8'b10001000;
    assign rom_data[2266]=8'b01100100;
    assign rom_data[2267]=8'b10001000;
    assign rom_data[2268]=8'b01100100;
    assign rom_data[2269]=8'b10000111;
    assign rom_data[2270]=8'b01100100;
    assign rom_data[2271]=8'b10000111;
    assign rom_data[2272]=8'b01100100;
    assign rom_data[2273]=8'b10000110;
    assign rom_data[2274]=8'b01100100;
    assign rom_data[2275]=8'b10000101;
    assign rom_data[2276]=8'b01100100;
    assign rom_data[2277]=8'b10000100;
    assign rom_data[2278]=8'b01100011;
    assign rom_data[2279]=8'b10000011;
    assign rom_data[2280]=8'b01100011;
    assign rom_data[2281]=8'b10000011;
    assign rom_data[2282]=8'b01100011;
    assign rom_data[2283]=8'b10000010;
    assign rom_data[2284]=8'b01100011;
    assign rom_data[2285]=8'b10000001;
    assign rom_data[2286]=8'b01100011;
    assign rom_data[2287]=8'b10000000;
    assign rom_data[2288]=8'b01100011;
    assign rom_data[2289]=8'b01111110;
    assign rom_data[2290]=8'b01100011;
    assign rom_data[2291]=8'b01111101;
    assign rom_data[2292]=8'b01100011;
    assign rom_data[2293]=8'b01111100;
    assign rom_data[2294]=8'b01100011;
    assign rom_data[2295]=8'b01111011;
    assign rom_data[2296]=8'b01100010;
    assign rom_data[2297]=8'b01111010;
    assign rom_data[2298]=8'b01100010;
    assign rom_data[2299]=8'b01111001;
    assign rom_data[2300]=8'b01100010;
    assign rom_data[2301]=8'b01110111;
    assign rom_data[2302]=8'b01100010;
    assign rom_data[2303]=8'b01110110;
    assign rom_data[2304]=8'b01100010;
    assign rom_data[2305]=8'b01110101;
    assign rom_data[2306]=8'b01100010;
    assign rom_data[2307]=8'b01110100;
    assign rom_data[2308]=8'b01100010;
    assign rom_data[2309]=8'b01110010;
    assign rom_data[2310]=8'b01100010;
    assign rom_data[2311]=8'b01110001;
    assign rom_data[2312]=8'b01100010;
    assign rom_data[2313]=8'b01110000;
    assign rom_data[2314]=8'b01100001;
    assign rom_data[2315]=8'b01101110;
    assign rom_data[2316]=8'b01100001;
    assign rom_data[2317]=8'b01101101;
    assign rom_data[2318]=8'b01100001;
    assign rom_data[2319]=8'b01101100;
    assign rom_data[2320]=8'b01100001;
    assign rom_data[2321]=8'b01101010;
    assign rom_data[2322]=8'b01100001;
    assign rom_data[2323]=8'b01101001;
    assign rom_data[2324]=8'b01100001;
    assign rom_data[2325]=8'b01100111;
    assign rom_data[2326]=8'b01100001;
    assign rom_data[2327]=8'b01100110;
    assign rom_data[2328]=8'b01100001;
    assign rom_data[2329]=8'b01100101;
    assign rom_data[2330]=8'b01100001;
    assign rom_data[2331]=8'b01100011;
    assign rom_data[2332]=8'b01100001;
    assign rom_data[2333]=8'b01100010;
    assign rom_data[2334]=8'b01100000;
    assign rom_data[2335]=8'b01100001;
    assign rom_data[2336]=8'b01100000;
    assign rom_data[2337]=8'b01011111;
    assign rom_data[2338]=8'b01100000;
    assign rom_data[2339]=8'b01011110;
    assign rom_data[2340]=8'b01100000;
    assign rom_data[2341]=8'b01011100;
    assign rom_data[2342]=8'b01100000;
    assign rom_data[2343]=8'b01011011;
    assign rom_data[2344]=8'b01100000;
    assign rom_data[2345]=8'b01011001;
    assign rom_data[2346]=8'b01100000;
    assign rom_data[2347]=8'b01011000;
    assign rom_data[2348]=8'b01100000;
    assign rom_data[2349]=8'b01010111;
    assign rom_data[2350]=8'b01100000;
    assign rom_data[2351]=8'b01010101;
    assign rom_data[2352]=8'b01100000;
    assign rom_data[2353]=8'b01010100;
    assign rom_data[2354]=8'b01011111;
    assign rom_data[2355]=8'b01010010;
    assign rom_data[2356]=8'b01011111;
    assign rom_data[2357]=8'b01010001;
    assign rom_data[2358]=8'b01011111;
    assign rom_data[2359]=8'b01010000;
    assign rom_data[2360]=8'b01011111;
    assign rom_data[2361]=8'b01001110;
    assign rom_data[2362]=8'b01011111;
    assign rom_data[2363]=8'b01001101;
    assign rom_data[2364]=8'b01011111;
    assign rom_data[2365]=8'b01001100;
    assign rom_data[2366]=8'b01011111;
    assign rom_data[2367]=8'b01001010;
    assign rom_data[2368]=8'b01011111;
    assign rom_data[2369]=8'b01001001;
    assign rom_data[2370]=8'b01011111;
    assign rom_data[2371]=8'b01001000;
    assign rom_data[2372]=8'b01011111;
    assign rom_data[2373]=8'b01000110;
    assign rom_data[2374]=8'b01011110;
    assign rom_data[2375]=8'b01000101;
    assign rom_data[2376]=8'b01011110;
    assign rom_data[2377]=8'b01000100;
    assign rom_data[2378]=8'b01011110;
    assign rom_data[2379]=8'b01000010;
    assign rom_data[2380]=8'b01011110;
    assign rom_data[2381]=8'b01000001;
    assign rom_data[2382]=8'b01011110;
    assign rom_data[2383]=8'b01000000;
    assign rom_data[2384]=8'b01011110;
    assign rom_data[2385]=8'b00111111;
    assign rom_data[2386]=8'b01011110;
    assign rom_data[2387]=8'b00111101;
    assign rom_data[2388]=8'b01011110;
    assign rom_data[2389]=8'b00111100;
    assign rom_data[2390]=8'b01011110;
    assign rom_data[2391]=8'b00111011;
    assign rom_data[2392]=8'b01011101;
    assign rom_data[2393]=8'b00111010;
    assign rom_data[2394]=8'b01011101;
    assign rom_data[2395]=8'b00111001;
    assign rom_data[2396]=8'b01011101;
    assign rom_data[2397]=8'b00111000;
    assign rom_data[2398]=8'b01011101;
    assign rom_data[2399]=8'b00110110;
    assign rom_data[2400]=8'b01011101;
    assign rom_data[2401]=8'b00110101;
    assign rom_data[2402]=8'b01011101;
    assign rom_data[2403]=8'b00110100;
    assign rom_data[2404]=8'b01011101;
    assign rom_data[2405]=8'b00110011;
    assign rom_data[2406]=8'b01011101;
    assign rom_data[2407]=8'b00110011;
    assign rom_data[2408]=8'b01011100;
    assign rom_data[2409]=8'b00110010;
    assign rom_data[2410]=8'b01011100;
    assign rom_data[2411]=8'b00110001;
    assign rom_data[2412]=8'b01011100;
    assign rom_data[2413]=8'b00110000;
    assign rom_data[2414]=8'b01011100;
    assign rom_data[2415]=8'b00101111;
    assign rom_data[2416]=8'b01011100;
    assign rom_data[2417]=8'b00101111;
    assign rom_data[2418]=8'b01011100;
    assign rom_data[2419]=8'b00101110;
    assign rom_data[2420]=8'b01011100;
    assign rom_data[2421]=8'b00101110;
    assign rom_data[2422]=8'b01011011;
    assign rom_data[2423]=8'b00101101;
    assign rom_data[2424]=8'b01011011;
    assign rom_data[2425]=8'b00101101;
    assign rom_data[2426]=8'b01011011;
    assign rom_data[2427]=8'b00101100;
    assign rom_data[2428]=8'b01011011;
    assign rom_data[2429]=8'b00101100;
    assign rom_data[2430]=8'b01011011;
    assign rom_data[2431]=8'b00101100;
    assign rom_data[2432]=8'b01011011;
    assign rom_data[2433]=8'b00101100;
    assign rom_data[2434]=8'b01011011;
    assign rom_data[2435]=8'b00101100;
    assign rom_data[2436]=8'b01011011;
    assign rom_data[2437]=8'b00101100;
    assign rom_data[2438]=8'b01011010;
    assign rom_data[2439]=8'b00101100;
    assign rom_data[2440]=8'b01011010;
    assign rom_data[2441]=8'b00101101;
    assign rom_data[2442]=8'b01011010;
    assign rom_data[2443]=8'b00101101;
    assign rom_data[2444]=8'b01011010;
    assign rom_data[2445]=8'b00101101;
    assign rom_data[2446]=8'b01011010;
    assign rom_data[2447]=8'b00101110;
    assign rom_data[2448]=8'b01011010;
    assign rom_data[2449]=8'b00101111;
    assign rom_data[2450]=8'b01011010;
    assign rom_data[2451]=8'b00101111;
    assign rom_data[2452]=8'b01011001;
    assign rom_data[2453]=8'b00110000;
    assign rom_data[2454]=8'b01011001;
    assign rom_data[2455]=8'b00110001;
    assign rom_data[2456]=8'b01011001;
    assign rom_data[2457]=8'b00110001;
    assign rom_data[2458]=8'b01011001;
    assign rom_data[2459]=8'b00110010;
    assign rom_data[2460]=8'b01011001;
    assign rom_data[2461]=8'b00110011;
    assign rom_data[2462]=8'b01011001;
    assign rom_data[2463]=8'b00110100;
    assign rom_data[2464]=8'b01011001;
    assign rom_data[2465]=8'b00110101;
    assign rom_data[2466]=8'b01011001;
    assign rom_data[2467]=8'b00110110;
    assign rom_data[2468]=8'b01011000;
    assign rom_data[2469]=8'b00110111;
    assign rom_data[2470]=8'b01011000;
    assign rom_data[2471]=8'b00111000;
    assign rom_data[2472]=8'b01011000;
    assign rom_data[2473]=8'b00111010;
    assign rom_data[2474]=8'b01011000;
    assign rom_data[2475]=8'b00111011;
    assign rom_data[2476]=8'b01011000;
    assign rom_data[2477]=8'b00111100;
    assign rom_data[2478]=8'b01011000;
    assign rom_data[2479]=8'b00111101;
    assign rom_data[2480]=8'b01011000;
    assign rom_data[2481]=8'b00111110;
    assign rom_data[2482]=8'b01011000;
    assign rom_data[2483]=8'b01000000;
    assign rom_data[2484]=8'b01011000;
    assign rom_data[2485]=8'b01000001;
    assign rom_data[2486]=8'b01010111;
    assign rom_data[2487]=8'b01000010;
    assign rom_data[2488]=8'b01010111;
    assign rom_data[2489]=8'b01000100;
    assign rom_data[2490]=8'b01010111;
    assign rom_data[2491]=8'b01000101;
    assign rom_data[2492]=8'b01010111;
    assign rom_data[2493]=8'b01000110;
    assign rom_data[2494]=8'b01010111;
    assign rom_data[2495]=8'b01000111;
    assign rom_data[2496]=8'b01010111;
    assign rom_data[2497]=8'b01001001;
    assign rom_data[2498]=8'b01010111;
    assign rom_data[2499]=8'b01001010;
    assign rom_data[2500]=8'b01010111;
    assign rom_data[2501]=8'b01001100;
    assign rom_data[2502]=8'b01010111;
    assign rom_data[2503]=8'b01001101;
    assign rom_data[2504]=8'b01010111;
    assign rom_data[2505]=8'b01001110;
    assign rom_data[2506]=8'b01010110;
    assign rom_data[2507]=8'b01010000;
    assign rom_data[2508]=8'b01010110;
    assign rom_data[2509]=8'b01010001;
    assign rom_data[2510]=8'b01010110;
    assign rom_data[2511]=8'b01010010;
    assign rom_data[2512]=8'b01010110;
    assign rom_data[2513]=8'b01010100;
    assign rom_data[2514]=8'b01010110;
    assign rom_data[2515]=8'b01010101;
    assign rom_data[2516]=8'b01010110;
    assign rom_data[2517]=8'b01010111;
    assign rom_data[2518]=8'b01010110;
    assign rom_data[2519]=8'b01011000;
    assign rom_data[2520]=8'b01010110;
    assign rom_data[2521]=8'b01011010;
    assign rom_data[2522]=8'b01010110;
    assign rom_data[2523]=8'b01011011;
    assign rom_data[2524]=8'b01010110;
    assign rom_data[2525]=8'b01011100;
    assign rom_data[2526]=8'b01010101;
    assign rom_data[2527]=8'b01011110;
    assign rom_data[2528]=8'b01010101;
    assign rom_data[2529]=8'b01011111;
    assign rom_data[2530]=8'b01010101;
    assign rom_data[2531]=8'b01100001;
    assign rom_data[2532]=8'b01010101;
    assign rom_data[2533]=8'b01100010;
    assign rom_data[2534]=8'b01010101;
    assign rom_data[2535]=8'b01100011;
    assign rom_data[2536]=8'b01010101;
    assign rom_data[2537]=8'b01100101;
    assign rom_data[2538]=8'b01010101;
    assign rom_data[2539]=8'b01100110;
    assign rom_data[2540]=8'b01010101;
    assign rom_data[2541]=8'b01100111;
    assign rom_data[2542]=8'b01010101;
    assign rom_data[2543]=8'b01101001;
    assign rom_data[2544]=8'b01010101;
    assign rom_data[2545]=8'b01101010;
    assign rom_data[2546]=8'b01010100;
    assign rom_data[2547]=8'b01101100;
    assign rom_data[2548]=8'b01010100;
    assign rom_data[2549]=8'b01101101;
    assign rom_data[2550]=8'b01010100;
    assign rom_data[2551]=8'b01101110;
    assign rom_data[2552]=8'b01010100;
    assign rom_data[2553]=8'b01110000;
    assign rom_data[2554]=8'b01010100;
    assign rom_data[2555]=8'b01110001;
    assign rom_data[2556]=8'b01010100;
    assign rom_data[2557]=8'b01110010;
    assign rom_data[2558]=8'b01010100;
    assign rom_data[2559]=8'b01110100;
    assign rom_data[2560]=8'b01010100;
    assign rom_data[2561]=8'b01110101;
    assign rom_data[2562]=8'b01010100;
    assign rom_data[2563]=8'b01110110;
    assign rom_data[2564]=8'b01010011;
    assign rom_data[2565]=8'b01110111;
    assign rom_data[2566]=8'b01010011;
    assign rom_data[2567]=8'b01111001;
    assign rom_data[2568]=8'b01010011;
    assign rom_data[2569]=8'b01111010;
    assign rom_data[2570]=8'b01010011;
    assign rom_data[2571]=8'b01111011;
    assign rom_data[2572]=8'b01010011;
    assign rom_data[2573]=8'b01111100;
    assign rom_data[2574]=8'b01010011;
    assign rom_data[2575]=8'b01111101;
    assign rom_data[2576]=8'b01010011;
    assign rom_data[2577]=8'b01111110;
    assign rom_data[2578]=8'b01010011;
    assign rom_data[2579]=8'b01111111;
    assign rom_data[2580]=8'b01010011;
    assign rom_data[2581]=8'b10000000;
    assign rom_data[2582]=8'b01010010;
    assign rom_data[2583]=8'b10000001;
    assign rom_data[2584]=8'b01010010;
    assign rom_data[2585]=8'b10000010;
    assign rom_data[2586]=8'b01010010;
    assign rom_data[2587]=8'b10000011;
    assign rom_data[2588]=8'b01010010;
    assign rom_data[2589]=8'b10000100;
    assign rom_data[2590]=8'b01010010;
    assign rom_data[2591]=8'b10000101;
    assign rom_data[2592]=8'b01010010;
    assign rom_data[2593]=8'b10000110;
    assign rom_data[2594]=8'b01010010;
    assign rom_data[2595]=8'b10000110;
    assign rom_data[2596]=8'b01010001;
    assign rom_data[2597]=8'b10000111;
    assign rom_data[2598]=8'b01010001;
    assign rom_data[2599]=8'b10001000;
    assign rom_data[2600]=8'b01010001;
    assign rom_data[2601]=8'b10001000;
    assign rom_data[2602]=8'b01010001;
    assign rom_data[2603]=8'b10001001;
    assign rom_data[2604]=8'b01010001;
    assign rom_data[2605]=8'b10001001;
    assign rom_data[2606]=8'b01010001;
    assign rom_data[2607]=8'b10001001;
    assign rom_data[2608]=8'b01010001;
    assign rom_data[2609]=8'b10001010;
    assign rom_data[2610]=8'b01010001;
    assign rom_data[2611]=8'b10001010;
    assign rom_data[2612]=8'b01010000;
    assign rom_data[2613]=8'b10001010;
    assign rom_data[2614]=8'b01010000;
    assign rom_data[2615]=8'b10001010;
    assign rom_data[2616]=8'b01010000;
    assign rom_data[2617]=8'b10001010;
    assign rom_data[2618]=8'b01010000;
    assign rom_data[2619]=8'b10001001;
    assign rom_data[2620]=8'b01010000;
    assign rom_data[2621]=8'b10001001;
    assign rom_data[2622]=8'b01010000;
    assign rom_data[2623]=8'b10001001;
    assign rom_data[2624]=8'b01010000;
    assign rom_data[2625]=8'b10001000;
    assign rom_data[2626]=8'b01001111;
    assign rom_data[2627]=8'b10001000;
    assign rom_data[2628]=8'b01001111;
    assign rom_data[2629]=8'b10000111;
    assign rom_data[2630]=8'b01001111;
    assign rom_data[2631]=8'b10000111;
    assign rom_data[2632]=8'b01001111;
    assign rom_data[2633]=8'b10000110;
    assign rom_data[2634]=8'b01001111;
    assign rom_data[2635]=8'b10000101;
    assign rom_data[2636]=8'b01001111;
    assign rom_data[2637]=8'b10000100;
    assign rom_data[2638]=8'b01001111;
    assign rom_data[2639]=8'b10000011;
    assign rom_data[2640]=8'b01001111;
    assign rom_data[2641]=8'b10000011;
    assign rom_data[2642]=8'b01001110;
    assign rom_data[2643]=8'b10000010;
    assign rom_data[2644]=8'b01001110;
    assign rom_data[2645]=8'b10000001;
    assign rom_data[2646]=8'b01001110;
    assign rom_data[2647]=8'b10000000;
    assign rom_data[2648]=8'b01001110;
    assign rom_data[2649]=8'b01111110;
    assign rom_data[2650]=8'b01001110;
    assign rom_data[2651]=8'b01111101;
    assign rom_data[2652]=8'b01001110;
    assign rom_data[2653]=8'b01111100;
    assign rom_data[2654]=8'b01001110;
    assign rom_data[2655]=8'b01111011;
    assign rom_data[2656]=8'b01001110;
    assign rom_data[2657]=8'b01111010;
    assign rom_data[2658]=8'b01001101;
    assign rom_data[2659]=8'b01111001;
    assign rom_data[2660]=8'b01001101;
    assign rom_data[2661]=8'b01110111;
    assign rom_data[2662]=8'b01001101;
    assign rom_data[2663]=8'b01110110;
    assign rom_data[2664]=8'b01001101;
    assign rom_data[2665]=8'b01110101;
    assign rom_data[2666]=8'b01001101;
    assign rom_data[2667]=8'b01110100;
    assign rom_data[2668]=8'b01001101;
    assign rom_data[2669]=8'b01110010;
    assign rom_data[2670]=8'b01001101;
    assign rom_data[2671]=8'b01110001;
    assign rom_data[2672]=8'b01001101;
    assign rom_data[2673]=8'b01110000;
    assign rom_data[2674]=8'b01001101;
    assign rom_data[2675]=8'b01101110;
    assign rom_data[2676]=8'b01001101;
    assign rom_data[2677]=8'b01101101;
    assign rom_data[2678]=8'b01001100;
    assign rom_data[2679]=8'b01101100;
    assign rom_data[2680]=8'b01001100;
    assign rom_data[2681]=8'b01101010;
    assign rom_data[2682]=8'b01001100;
    assign rom_data[2683]=8'b01101001;
    assign rom_data[2684]=8'b01001100;
    assign rom_data[2685]=8'b01100111;
    assign rom_data[2686]=8'b01001100;
    assign rom_data[2687]=8'b01100110;
    assign rom_data[2688]=8'b01001100;
    assign rom_data[2689]=8'b01100101;
    assign rom_data[2690]=8'b01001100;
    assign rom_data[2691]=8'b01100011;
    assign rom_data[2692]=8'b01001100;
    assign rom_data[2693]=8'b01100010;
    assign rom_data[2694]=8'b01001100;
    assign rom_data[2695]=8'b01100001;
    assign rom_data[2696]=8'b01001100;
    assign rom_data[2697]=8'b01011111;
    assign rom_data[2698]=8'b01001011;
    assign rom_data[2699]=8'b01011110;
    assign rom_data[2700]=8'b01001011;
    assign rom_data[2701]=8'b01011100;
    assign rom_data[2702]=8'b01001011;
    assign rom_data[2703]=8'b01011011;
    assign rom_data[2704]=8'b01001011;
    assign rom_data[2705]=8'b01011001;
    assign rom_data[2706]=8'b01001011;
    assign rom_data[2707]=8'b01011000;
    assign rom_data[2708]=8'b01001011;
    assign rom_data[2709]=8'b01010111;
    assign rom_data[2710]=8'b01001011;
    assign rom_data[2711]=8'b01010101;
    assign rom_data[2712]=8'b01001011;
    assign rom_data[2713]=8'b01010100;
    assign rom_data[2714]=8'b01001011;
    assign rom_data[2715]=8'b01010010;
    assign rom_data[2716]=8'b01001011;
    assign rom_data[2717]=8'b01010001;
    assign rom_data[2718]=8'b01001010;
    assign rom_data[2719]=8'b01010000;
    assign rom_data[2720]=8'b01001010;
    assign rom_data[2721]=8'b01001110;
    assign rom_data[2722]=8'b01001010;
    assign rom_data[2723]=8'b01001101;
    assign rom_data[2724]=8'b01001010;
    assign rom_data[2725]=8'b01001100;
    assign rom_data[2726]=8'b01001010;
    assign rom_data[2727]=8'b01001010;
    assign rom_data[2728]=8'b01001010;
    assign rom_data[2729]=8'b01001001;
    assign rom_data[2730]=8'b01001010;
    assign rom_data[2731]=8'b01001000;
    assign rom_data[2732]=8'b01001010;
    assign rom_data[2733]=8'b01000110;
    assign rom_data[2734]=8'b01001010;
    assign rom_data[2735]=8'b01000101;
    assign rom_data[2736]=8'b01001001;
    assign rom_data[2737]=8'b01000100;
    assign rom_data[2738]=8'b01001001;
    assign rom_data[2739]=8'b01000010;
    assign rom_data[2740]=8'b01001001;
    assign rom_data[2741]=8'b01000001;
    assign rom_data[2742]=8'b01001001;
    assign rom_data[2743]=8'b01000000;
    assign rom_data[2744]=8'b01001001;
    assign rom_data[2745]=8'b00111111;
    assign rom_data[2746]=8'b01001001;
    assign rom_data[2747]=8'b00111101;
    assign rom_data[2748]=8'b01001001;
    assign rom_data[2749]=8'b00111100;
    assign rom_data[2750]=8'b01001001;
    assign rom_data[2751]=8'b00111011;
    assign rom_data[2752]=8'b01001001;
    assign rom_data[2753]=8'b00111010;
    assign rom_data[2754]=8'b01001000;
    assign rom_data[2755]=8'b00111001;
    assign rom_data[2756]=8'b01001000;
    assign rom_data[2757]=8'b00111000;
    assign rom_data[2758]=8'b01001000;
    assign rom_data[2759]=8'b00110110;
    assign rom_data[2760]=8'b01001000;
    assign rom_data[2761]=8'b00110101;
    assign rom_data[2762]=8'b01001000;
    assign rom_data[2763]=8'b00110100;
    assign rom_data[2764]=8'b01001000;
    assign rom_data[2765]=8'b00110011;
    assign rom_data[2766]=8'b01001000;
    assign rom_data[2767]=8'b00110011;
    assign rom_data[2768]=8'b01001000;
    assign rom_data[2769]=8'b00110010;
    assign rom_data[2770]=8'b01000111;
    assign rom_data[2771]=8'b00110001;
    assign rom_data[2772]=8'b01000111;
    assign rom_data[2773]=8'b00110000;
    assign rom_data[2774]=8'b01000111;
    assign rom_data[2775]=8'b00101111;
    assign rom_data[2776]=8'b01000111;
    assign rom_data[2777]=8'b00101111;
    assign rom_data[2778]=8'b01000111;
    assign rom_data[2779]=8'b00101110;
    assign rom_data[2780]=8'b01000111;
    assign rom_data[2781]=8'b00101110;
    assign rom_data[2782]=8'b01000111;
    assign rom_data[2783]=8'b00101101;
    assign rom_data[2784]=8'b01000111;
    assign rom_data[2785]=8'b00101101;
    assign rom_data[2786]=8'b01000110;
    assign rom_data[2787]=8'b00101100;
    assign rom_data[2788]=8'b01000110;
    assign rom_data[2789]=8'b00101100;
    assign rom_data[2790]=8'b01000110;
    assign rom_data[2791]=8'b00101100;
    assign rom_data[2792]=8'b01000110;
    assign rom_data[2793]=8'b00101100;
    assign rom_data[2794]=8'b01000110;
    assign rom_data[2795]=8'b00101100;
    assign rom_data[2796]=8'b01000110;
    assign rom_data[2797]=8'b00101100;
    assign rom_data[2798]=8'b01000110;
    assign rom_data[2799]=8'b00101100;
    assign rom_data[2800]=8'b01000101;
    assign rom_data[2801]=8'b00101101;
    assign rom_data[2802]=8'b01000101;
    assign rom_data[2803]=8'b00101101;
    assign rom_data[2804]=8'b01000101;
    assign rom_data[2805]=8'b00101101;
    assign rom_data[2806]=8'b01000101;
    assign rom_data[2807]=8'b00101110;
    assign rom_data[2808]=8'b01000101;
    assign rom_data[2809]=8'b00101111;
    assign rom_data[2810]=8'b01000101;
    assign rom_data[2811]=8'b00101111;
    assign rom_data[2812]=8'b01000101;
    assign rom_data[2813]=8'b00110000;
    assign rom_data[2814]=8'b01000100;
    assign rom_data[2815]=8'b00110001;
    assign rom_data[2816]=8'b01000100;
    assign rom_data[2817]=8'b00110001;
    assign rom_data[2818]=8'b01000100;
    assign rom_data[2819]=8'b00110010;
    assign rom_data[2820]=8'b01000100;
    assign rom_data[2821]=8'b00110011;
    assign rom_data[2822]=8'b01000100;
    assign rom_data[2823]=8'b00110100;
    assign rom_data[2824]=8'b01000100;
    assign rom_data[2825]=8'b00110101;
    assign rom_data[2826]=8'b01000100;
    assign rom_data[2827]=8'b00110110;
    assign rom_data[2828]=8'b01000100;
    assign rom_data[2829]=8'b00110111;
    assign rom_data[2830]=8'b01000011;
    assign rom_data[2831]=8'b00111000;
    assign rom_data[2832]=8'b01000011;
    assign rom_data[2833]=8'b00111010;
    assign rom_data[2834]=8'b01000011;
    assign rom_data[2835]=8'b00111011;
    assign rom_data[2836]=8'b01000011;
    assign rom_data[2837]=8'b00111100;
    assign rom_data[2838]=8'b01000011;
    assign rom_data[2839]=8'b00111101;
    assign rom_data[2840]=8'b01000011;
    assign rom_data[2841]=8'b00111110;
    assign rom_data[2842]=8'b01000011;
    assign rom_data[2843]=8'b01000000;
    assign rom_data[2844]=8'b01000011;
    assign rom_data[2845]=8'b01000001;
    assign rom_data[2846]=8'b01000011;
    assign rom_data[2847]=8'b01000010;
    assign rom_data[2848]=8'b01000011;
    assign rom_data[2849]=8'b01000100;
    assign rom_data[2850]=8'b01000010;
    assign rom_data[2851]=8'b01000101;
    assign rom_data[2852]=8'b01000010;
    assign rom_data[2853]=8'b01000110;
    assign rom_data[2854]=8'b01000010;
    assign rom_data[2855]=8'b01000111;
    assign rom_data[2856]=8'b01000010;
    assign rom_data[2857]=8'b01001001;
    assign rom_data[2858]=8'b01000010;
    assign rom_data[2859]=8'b01001010;
    assign rom_data[2860]=8'b01000010;
    assign rom_data[2861]=8'b01001100;
    assign rom_data[2862]=8'b01000010;
    assign rom_data[2863]=8'b01001101;
    assign rom_data[2864]=8'b01000010;
    assign rom_data[2865]=8'b01001110;
    assign rom_data[2866]=8'b01000010;
    assign rom_data[2867]=8'b01010000;
    assign rom_data[2868]=8'b01000001;
    assign rom_data[2869]=8'b01010001;
    assign rom_data[2870]=8'b01000001;
    assign rom_data[2871]=8'b01010010;
    assign rom_data[2872]=8'b01000001;
    assign rom_data[2873]=8'b01010100;
    assign rom_data[2874]=8'b01000001;
    assign rom_data[2875]=8'b01010101;
    assign rom_data[2876]=8'b01000001;
    assign rom_data[2877]=8'b01010111;
    assign rom_data[2878]=8'b01000001;
    assign rom_data[2879]=8'b01011000;
    assign rom_data[2880]=8'b01000001;
    assign rom_data[2881]=8'b01011010;
    assign rom_data[2882]=8'b01000001;
    assign rom_data[2883]=8'b01011011;
    assign rom_data[2884]=8'b01000001;
    assign rom_data[2885]=8'b01011100;
    assign rom_data[2886]=8'b01000001;
    assign rom_data[2887]=8'b01011110;
    assign rom_data[2888]=8'b01000000;
    assign rom_data[2889]=8'b01011111;
    assign rom_data[2890]=8'b01000000;
    assign rom_data[2891]=8'b01100001;
    assign rom_data[2892]=8'b01000000;
    assign rom_data[2893]=8'b01100010;
    assign rom_data[2894]=8'b01000000;
    assign rom_data[2895]=8'b01100011;
    assign rom_data[2896]=8'b01000000;
    assign rom_data[2897]=8'b01100101;
    assign rom_data[2898]=8'b01000000;
    assign rom_data[2899]=8'b01100110;
    assign rom_data[2900]=8'b01000000;
    assign rom_data[2901]=8'b01100111;
    assign rom_data[2902]=8'b01000000;
    assign rom_data[2903]=8'b01101001;
    assign rom_data[2904]=8'b01000000;
    assign rom_data[2905]=8'b01101010;
    assign rom_data[2906]=8'b01000000;
    assign rom_data[2907]=8'b01101100;
    assign rom_data[2908]=8'b00111111;
    assign rom_data[2909]=8'b01101101;
    assign rom_data[2910]=8'b00111111;
    assign rom_data[2911]=8'b01101110;
    assign rom_data[2912]=8'b00111111;
    assign rom_data[2913]=8'b01110000;
    assign rom_data[2914]=8'b00111111;
    assign rom_data[2915]=8'b01110001;
    assign rom_data[2916]=8'b00111111;
    assign rom_data[2917]=8'b01110010;
    assign rom_data[2918]=8'b00111111;
    assign rom_data[2919]=8'b01110100;
    assign rom_data[2920]=8'b00111111;
    assign rom_data[2921]=8'b01110101;
    assign rom_data[2922]=8'b00111111;
    assign rom_data[2923]=8'b01110110;
    assign rom_data[2924]=8'b00111111;
    assign rom_data[2925]=8'b01110111;
    assign rom_data[2926]=8'b00111110;
    assign rom_data[2927]=8'b01111001;
    assign rom_data[2928]=8'b00111110;
    assign rom_data[2929]=8'b01111010;
    assign rom_data[2930]=8'b00111110;
    assign rom_data[2931]=8'b01111011;
    assign rom_data[2932]=8'b00111110;
    assign rom_data[2933]=8'b01111100;
    assign rom_data[2934]=8'b00111110;
    assign rom_data[2935]=8'b01111101;
    assign rom_data[2936]=8'b00111110;
    assign rom_data[2937]=8'b01111110;
    assign rom_data[2938]=8'b00111110;
    assign rom_data[2939]=8'b01111111;
    assign rom_data[2940]=8'b00111110;
    assign rom_data[2941]=8'b10000000;
    assign rom_data[2942]=8'b00111110;
    assign rom_data[2943]=8'b10000001;
    assign rom_data[2944]=8'b00111101;
    assign rom_data[2945]=8'b10000010;
    assign rom_data[2946]=8'b00111101;
    assign rom_data[2947]=8'b10000011;
    assign rom_data[2948]=8'b00111101;
    assign rom_data[2949]=8'b10000100;
    assign rom_data[2950]=8'b00111101;
    assign rom_data[2951]=8'b10000101;
    assign rom_data[2952]=8'b00111101;
    assign rom_data[2953]=8'b10000110;
    assign rom_data[2954]=8'b00111101;
    assign rom_data[2955]=8'b10000110;
    assign rom_data[2956]=8'b00111101;
    assign rom_data[2957]=8'b10000111;
    assign rom_data[2958]=8'b00111100;
    assign rom_data[2959]=8'b10001000;
    assign rom_data[2960]=8'b00111100;
    assign rom_data[2961]=8'b10001000;
    assign rom_data[2962]=8'b00111100;
    assign rom_data[2963]=8'b10001001;
    assign rom_data[2964]=8'b00111100;
    assign rom_data[2965]=8'b10001001;
    assign rom_data[2966]=8'b00111100;
    assign rom_data[2967]=8'b10001001;
    assign rom_data[2968]=8'b00111100;
    assign rom_data[2969]=8'b10001010;
    assign rom_data[2970]=8'b00111100;
    assign rom_data[2971]=8'b10001010;
    assign rom_data[2972]=8'b00111100;
    assign rom_data[2973]=8'b10001010;
    assign rom_data[2974]=8'b00111011;
    assign rom_data[2975]=8'b10001010;
    assign rom_data[2976]=8'b00111011;
    assign rom_data[2977]=8'b10001010;
    assign rom_data[2978]=8'b00111011;
    assign rom_data[2979]=8'b10001001;
    assign rom_data[2980]=8'b00111011;
    assign rom_data[2981]=8'b10001001;
    assign rom_data[2982]=8'b00111011;
    assign rom_data[2983]=8'b10001001;
    assign rom_data[2984]=8'b00111011;
    assign rom_data[2985]=8'b10001000;
    assign rom_data[2986]=8'b00111011;
    assign rom_data[2987]=8'b10001000;
    assign rom_data[2988]=8'b00111010;
    assign rom_data[2989]=8'b10000111;
    assign rom_data[2990]=8'b00111010;
    assign rom_data[2991]=8'b10000111;
    assign rom_data[2992]=8'b00111010;
    assign rom_data[2993]=8'b10000110;
    assign rom_data[2994]=8'b00111010;
    assign rom_data[2995]=8'b10000101;
    assign rom_data[2996]=8'b00111010;
    assign rom_data[2997]=8'b10000100;
    assign rom_data[2998]=8'b00111010;
    assign rom_data[2999]=8'b10000011;
    assign rom_data[3000]=8'b00111010;
    assign rom_data[3001]=8'b10000011;
    assign rom_data[3002]=8'b00111010;
    assign rom_data[3003]=8'b10000010;
    assign rom_data[3004]=8'b00111001;
    assign rom_data[3005]=8'b10000001;
    assign rom_data[3006]=8'b00111001;
    assign rom_data[3007]=8'b10000000;
    assign rom_data[3008]=8'b00111001;
    assign rom_data[3009]=8'b01111110;
    assign rom_data[3010]=8'b00111001;
    assign rom_data[3011]=8'b01111101;
    assign rom_data[3012]=8'b00111001;
    assign rom_data[3013]=8'b01111100;
    assign rom_data[3014]=8'b00111001;
    assign rom_data[3015]=8'b01111011;
    assign rom_data[3016]=8'b00111001;
    assign rom_data[3017]=8'b01111010;
    assign rom_data[3018]=8'b00111001;
    assign rom_data[3019]=8'b01111001;
    assign rom_data[3020]=8'b00111001;
    assign rom_data[3021]=8'b01110111;
    assign rom_data[3022]=8'b00111000;
    assign rom_data[3023]=8'b01110110;
    assign rom_data[3024]=8'b00111000;
    assign rom_data[3025]=8'b01110101;
    assign rom_data[3026]=8'b00111000;
    assign rom_data[3027]=8'b01110100;
    assign rom_data[3028]=8'b00111000;
    assign rom_data[3029]=8'b01110010;
    assign rom_data[3030]=8'b00111000;
    assign rom_data[3031]=8'b01110001;
    assign rom_data[3032]=8'b00111000;
    assign rom_data[3033]=8'b01110000;
    assign rom_data[3034]=8'b00111000;
    assign rom_data[3035]=8'b01101110;
    assign rom_data[3036]=8'b00111000;
    assign rom_data[3037]=8'b01101101;
    assign rom_data[3038]=8'b00111000;
    assign rom_data[3039]=8'b01101100;
    assign rom_data[3040]=8'b00110111;
    assign rom_data[3041]=8'b01101010;
    assign rom_data[3042]=8'b00110111;
    assign rom_data[3043]=8'b01101001;
    assign rom_data[3044]=8'b00110111;
    assign rom_data[3045]=8'b01100111;
    assign rom_data[3046]=8'b00110111;
    assign rom_data[3047]=8'b01100110;
    assign rom_data[3048]=8'b00110111;
    assign rom_data[3049]=8'b01100101;
    assign rom_data[3050]=8'b00110111;
    assign rom_data[3051]=8'b01100011;
    assign rom_data[3052]=8'b00110111;
    assign rom_data[3053]=8'b01100010;
    assign rom_data[3054]=8'b00110111;
    assign rom_data[3055]=8'b01100001;
    assign rom_data[3056]=8'b00110111;
    assign rom_data[3057]=8'b01011111;
    assign rom_data[3058]=8'b00110111;
    assign rom_data[3059]=8'b01011110;
    assign rom_data[3060]=8'b00110110;
    assign rom_data[3061]=8'b01011100;
    assign rom_data[3062]=8'b00110110;
    assign rom_data[3063]=8'b01011011;
    assign rom_data[3064]=8'b00110110;
    assign rom_data[3065]=8'b01011001;
    assign rom_data[3066]=8'b00110110;
    assign rom_data[3067]=8'b01011000;
    assign rom_data[3068]=8'b00110110;
    assign rom_data[3069]=8'b01010111;
    assign rom_data[3070]=8'b00110110;
    assign rom_data[3071]=8'b01010101;
    assign rom_data[3072]=8'b00110110;
    assign rom_data[3073]=8'b01010100;
    assign rom_data[3074]=8'b00110110;
    assign rom_data[3075]=8'b01010010;
    assign rom_data[3076]=8'b00110110;
    assign rom_data[3077]=8'b01010001;
    assign rom_data[3078]=8'b00110110;
    assign rom_data[3079]=8'b01010000;
    assign rom_data[3080]=8'b00110101;
    assign rom_data[3081]=8'b01001110;
    assign rom_data[3082]=8'b00110101;
    assign rom_data[3083]=8'b01001101;
    assign rom_data[3084]=8'b00110101;
    assign rom_data[3085]=8'b01001100;
    assign rom_data[3086]=8'b00110101;
    assign rom_data[3087]=8'b01001010;
    assign rom_data[3088]=8'b00110101;
    assign rom_data[3089]=8'b01001001;
    assign rom_data[3090]=8'b00110101;
    assign rom_data[3091]=8'b01001000;
    assign rom_data[3092]=8'b00110101;
    assign rom_data[3093]=8'b01000110;
    assign rom_data[3094]=8'b00110101;
    assign rom_data[3095]=8'b01000101;
    assign rom_data[3096]=8'b00110101;
    assign rom_data[3097]=8'b01000100;
    assign rom_data[3098]=8'b00110101;
    assign rom_data[3099]=8'b01000010;
    assign rom_data[3100]=8'b00110100;
    assign rom_data[3101]=8'b01000001;
    assign rom_data[3102]=8'b00110100;
    assign rom_data[3103]=8'b01000000;
    assign rom_data[3104]=8'b00110100;
    assign rom_data[3105]=8'b00111111;
    assign rom_data[3106]=8'b00110100;
    assign rom_data[3107]=8'b00111101;
    assign rom_data[3108]=8'b00110100;
    assign rom_data[3109]=8'b00111100;
    assign rom_data[3110]=8'b00110100;
    assign rom_data[3111]=8'b00111011;
    assign rom_data[3112]=8'b00110100;
    assign rom_data[3113]=8'b00111010;
    assign rom_data[3114]=8'b00110100;
    assign rom_data[3115]=8'b00111001;
    assign rom_data[3116]=8'b00110011;
    assign rom_data[3117]=8'b00111000;
    assign rom_data[3118]=8'b00110011;
    assign rom_data[3119]=8'b00110110;
    assign rom_data[3120]=8'b00110011;
    assign rom_data[3121]=8'b00110101;
    assign rom_data[3122]=8'b00110011;
    assign rom_data[3123]=8'b00110100;
    assign rom_data[3124]=8'b00110011;
    assign rom_data[3125]=8'b00110011;
    assign rom_data[3126]=8'b00110011;
    assign rom_data[3127]=8'b00110011;
    assign rom_data[3128]=8'b00110011;
    assign rom_data[3129]=8'b00110010;
    assign rom_data[3130]=8'b00110011;
    assign rom_data[3131]=8'b00110001;
    assign rom_data[3132]=8'b00110010;
    assign rom_data[3133]=8'b00110000;
    assign rom_data[3134]=8'b00110010;
    assign rom_data[3135]=8'b00101111;
    assign rom_data[3136]=8'b00110010;
    assign rom_data[3137]=8'b00101111;
    assign rom_data[3138]=8'b00110010;
    assign rom_data[3139]=8'b00101110;
    assign rom_data[3140]=8'b00110010;
    assign rom_data[3141]=8'b00101110;
    assign rom_data[3142]=8'b00110010;
    assign rom_data[3143]=8'b00101101;
    assign rom_data[3144]=8'b00110010;
    assign rom_data[3145]=8'b00101101;
    assign rom_data[3146]=8'b00110010;
    assign rom_data[3147]=8'b00101100;
    assign rom_data[3148]=8'b00110001;
    assign rom_data[3149]=8'b00101100;
    assign rom_data[3150]=8'b00110001;
    assign rom_data[3151]=8'b00101100;
    assign rom_data[3152]=8'b00110001;
    assign rom_data[3153]=8'b00101100;
    assign rom_data[3154]=8'b00110001;
    assign rom_data[3155]=8'b00101100;
    assign rom_data[3156]=8'b00110001;
    assign rom_data[3157]=8'b00101100;
    assign rom_data[3158]=8'b00110001;
    assign rom_data[3159]=8'b00101100;
    assign rom_data[3160]=8'b00110001;
    assign rom_data[3161]=8'b00101101;
    assign rom_data[3162]=8'b00110000;
    assign rom_data[3163]=8'b00101101;
    assign rom_data[3164]=8'b00110000;
    assign rom_data[3165]=8'b00101101;
    assign rom_data[3166]=8'b00110000;
    assign rom_data[3167]=8'b00101110;
    assign rom_data[3168]=8'b00110000;
    assign rom_data[3169]=8'b00101111;
    assign rom_data[3170]=8'b00110000;
    assign rom_data[3171]=8'b00101111;
    assign rom_data[3172]=8'b00110000;
    assign rom_data[3173]=8'b00110000;
    assign rom_data[3174]=8'b00110000;
    assign rom_data[3175]=8'b00110001;
    assign rom_data[3176]=8'b00110000;
    assign rom_data[3177]=8'b00110001;
    assign rom_data[3178]=8'b00110000;
    assign rom_data[3179]=8'b00110010;
    assign rom_data[3180]=8'b00101111;
    assign rom_data[3181]=8'b00110011;
    assign rom_data[3182]=8'b00101111;
    assign rom_data[3183]=8'b00110100;
    assign rom_data[3184]=8'b00101111;
    assign rom_data[3185]=8'b00110101;
    assign rom_data[3186]=8'b00101111;
    assign rom_data[3187]=8'b00110110;
    assign rom_data[3188]=8'b00101111;
    assign rom_data[3189]=8'b00110111;
    assign rom_data[3190]=8'b00101111;
    assign rom_data[3191]=8'b00111000;
    assign rom_data[3192]=8'b00101111;
    assign rom_data[3193]=8'b00111010;
    assign rom_data[3194]=8'b00101111;
    assign rom_data[3195]=8'b00111011;
    assign rom_data[3196]=8'b00101111;
    assign rom_data[3197]=8'b00111100;
    assign rom_data[3198]=8'b00101110;
    assign rom_data[3199]=8'b00111101;
    assign rom_data[3200]=8'b00101110;
    assign rom_data[3201]=8'b00111110;
    assign rom_data[3202]=8'b00101110;
    assign rom_data[3203]=8'b01000000;
    assign rom_data[3204]=8'b00101110;
    assign rom_data[3205]=8'b01000001;
    assign rom_data[3206]=8'b00101110;
    assign rom_data[3207]=8'b01000010;
    assign rom_data[3208]=8'b00101110;
    assign rom_data[3209]=8'b01000100;
    assign rom_data[3210]=8'b00101110;
    assign rom_data[3211]=8'b01000101;
    assign rom_data[3212]=8'b00101110;
    assign rom_data[3213]=8'b01000110;
    assign rom_data[3214]=8'b00101110;
    assign rom_data[3215]=8'b01001000;
    assign rom_data[3216]=8'b00101110;
    assign rom_data[3217]=8'b01001001;
    assign rom_data[3218]=8'b00101110;
    assign rom_data[3219]=8'b01001010;
    assign rom_data[3220]=8'b00101110;
    assign rom_data[3221]=8'b01001100;
    assign rom_data[3222]=8'b00101110;
    assign rom_data[3223]=8'b01001101;
    assign rom_data[3224]=8'b00101110;
    assign rom_data[3225]=8'b01001110;
    assign rom_data[3226]=8'b00101101;
    assign rom_data[3227]=8'b01010000;
    assign rom_data[3228]=8'b00101101;
    assign rom_data[3229]=8'b01010001;
    assign rom_data[3230]=8'b00101101;
    assign rom_data[3231]=8'b01010010;
    assign rom_data[3232]=8'b00101101;
    assign rom_data[3233]=8'b01010100;
    assign rom_data[3234]=8'b00101101;
    assign rom_data[3235]=8'b01010101;
    assign rom_data[3236]=8'b00101101;
    assign rom_data[3237]=8'b01010111;
    assign rom_data[3238]=8'b00101101;
    assign rom_data[3239]=8'b01011000;
    assign rom_data[3240]=8'b00101101;
    assign rom_data[3241]=8'b01011010;


reg [23:0] f1_data_d, f1_data_q;
wire[13:0] f1_addrs;
reg [15:0] f1_antidata;

reg [23:0] f2_data_d, f2_data_q;
wire[13:0] f2_addrs;
reg [15:0] f2_antidata;

reg [23:0] f3_data_d, f3_data_q;
wire[13:0] f3_addrs;
reg [15:0] f3_antidata;

reg [23:0] f4_data_d, f4_data_q;
wire[13:0] f4_addrs;
reg [15:0] f4_antidata;

reg [23:0] f5_data_d, f5_data_q;
wire[13:0] f5_addrs;
reg [15:0] f5_antidata;

reg [23:0] f6_data_d, f6_data_q;
wire[13:0] f6_addrs;
reg [15:0] f6_antidata;

reg done;

reg [4:0] home_step=5'd30;
reg [15:0] home_bias=16'd23250;

reg [15:0] f1_CH_A_d, f1_CH_A_q;
reg [15:0] f1_CH_B_d, f1_CH_B_q;
reg [15:0] f1_CH_C_d, f1_CH_C_q;
reg [15:0] f1_CH_D_d, f1_CH_D_q;

reg [15:0] f2_CH_A_d, f2_CH_A_q;
reg [15:0] f2_CH_B_d, f2_CH_B_q;
reg [15:0] f2_CH_C_d, f2_CH_C_q;
reg [15:0] f2_CH_D_d, f2_CH_D_q;

reg [15:0] f3_CH_A_d, f3_CH_A_q;
reg [15:0] f3_CH_B_d, f3_CH_B_q;
reg [15:0] f3_CH_C_d, f3_CH_C_q;
reg [15:0] f3_CH_D_d, f3_CH_D_q;

reg [15:0] f4_CH_A_d, f4_CH_A_q;
reg [15:0] f4_CH_B_d, f4_CH_B_q;
reg [15:0] f4_CH_C_d, f4_CH_C_q;
reg [15:0] f4_CH_D_d, f4_CH_D_q;

reg [15:0] f5_CH_A_d, f5_CH_A_q;
reg [15:0] f5_CH_B_d, f5_CH_B_q;
reg [15:0] f5_CH_C_d, f5_CH_C_q;
reg [15:0] f5_CH_D_d, f5_CH_D_q;

reg [15:0] f6_CH_A_d, f6_CH_A_q;
reg [15:0] f6_CH_B_d, f6_CH_B_q;
reg [15:0] f6_CH_C_d, f6_CH_C_q;
reg [15:0] f6_CH_D_d, f6_CH_D_q;

assign f1_data = f1_data_q;
assign f2_data = f2_data_q;
assign f3_data = f3_data_q;
assign f4_data = f4_data_q;
assign f5_data = f5_data_q;
assign f6_data = f6_data_q;

assign f1_addrs = f1_addr[15:2];

assign f2_addrs = f2_addr[15:2];
assign f3_addrs = f3_addr[15:2];
assign f4_addrs = f4_addr[15:2];
assign f5_addrs = f5_addr[15:2];
assign f6_addrs = f6_addr[15:2];

always @(*) begin
    f1_CH_A_d=f1_CH_A_q;
    f1_CH_B_d=f1_CH_B_q;
    f1_CH_C_d=f1_CH_C_q;
    f1_CH_D_d=f1_CH_D_q;

    f2_CH_A_d=f2_CH_A_q;
    f2_CH_B_d=f2_CH_B_q;
    f2_CH_C_d=f2_CH_C_q;
    f2_CH_D_d=f2_CH_D_q;
    
    f3_CH_A_d=f3_CH_A_q;
    f3_CH_B_d=f3_CH_B_q;
    f3_CH_C_d=f3_CH_C_q;
    f3_CH_D_d=f3_CH_D_q;
    
    f4_CH_A_d=f4_CH_A_q;
    f4_CH_B_d=f4_CH_B_q;
    f4_CH_C_d=f4_CH_C_q;
    f4_CH_D_d=f4_CH_D_q;
    
    f5_CH_A_d=f5_CH_A_q;
    f5_CH_B_d=f5_CH_B_q;
    f5_CH_C_d=f5_CH_C_q;
    f5_CH_D_d=f5_CH_D_q;
    
    f6_CH_A_d=f6_CH_A_q;
    f6_CH_B_d=f6_CH_B_q;
    f6_CH_C_d=f6_CH_C_q;
    f6_CH_D_d=f6_CH_D_q;


    if (go_home==1'b1) begin
        // F1
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f1_CH_A_q>home_bias) begin
                    f1_CH_A_d=f1_CH_A_q-home_step;
                end else if (f1_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_A_d=f1_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f1_CH_C_q>home_bias) begin
                    f1_CH_C_d=f1_CH_C_q-home_step;
                end else if (f1_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_C_d=f1_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f1_CH_B_q>home_bias) begin
                    f1_CH_B_d=f1_CH_B_q-home_step;
                end else if (f1_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_B_d=f1_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f1_CH_D_q>home_bias) begin
                    f1_CH_D_d=f1_CH_D_q-home_step;
                end else if (f1_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f1_CH_D_d=f1_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f2_CH_A_q>home_bias) begin
                    f2_CH_A_d=f2_CH_A_q-home_step;
                end else if (f2_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_A_d=f2_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f2_CH_C_q>home_bias) begin
                    f2_CH_C_d=f2_CH_C_q-home_step;
                end else if (f2_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_C_d=f2_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f2_CH_B_q>home_bias) begin
                    f2_CH_B_d=f2_CH_B_q-home_step;
                end else if (f2_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_B_d=f2_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f2_CH_D_q>home_bias) begin
                    f2_CH_D_d=f2_CH_D_q-home_step;
                end else if (f2_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f2_CH_D_d=f2_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F3
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f3_CH_A_q>home_bias) begin
                    f3_CH_A_d=f3_CH_A_q-home_step;
                end else if (f3_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_A_d=f3_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f3_CH_C_q>home_bias) begin
                    f3_CH_C_d=f3_CH_C_q-home_step;
                end else if (f3_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_C_d=f3_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f3_CH_B_q>home_bias) begin
                    f3_CH_B_d=f3_CH_B_q-home_step;
                end else if (f3_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_B_d=f3_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f3_CH_D_q>home_bias) begin
                    f3_CH_D_d=f3_CH_D_q-home_step;
                end else if (f3_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f3_CH_D_d=f3_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F4
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f4_CH_A_q>home_bias) begin
                    f4_CH_A_d=f4_CH_A_q-home_step;
                end else if (f4_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_A_d=f4_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f4_CH_C_q>home_bias) begin
                    f4_CH_C_d=f4_CH_C_q-home_step;
                end else if (f4_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_C_d=f4_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f4_CH_B_q>home_bias) begin
                    f4_CH_B_d=f4_CH_B_q-home_step;
                end else if (f4_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_B_d=f4_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f4_CH_D_q>home_bias) begin
                    f4_CH_D_d=f4_CH_D_q-home_step;
                end else if (f4_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f4_CH_D_d=f4_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F5
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f5_CH_A_q>home_bias) begin
                    f5_CH_A_d=f5_CH_A_q-home_step;
                end else if (f5_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_A_d=f5_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f5_CH_C_q>home_bias) begin
                    f5_CH_C_d=f5_CH_C_q-home_step;
                end else if (f5_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_C_d=f5_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f5_CH_B_q>home_bias) begin
                    f5_CH_B_d=f5_CH_B_q-home_step;
                end else if (f5_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_B_d=f5_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f5_CH_D_q>home_bias) begin
                    f5_CH_D_d=f5_CH_D_q-home_step;
                end else if (f5_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f5_CH_D_d=f5_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
        // F6
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                if (f6_CH_A_q>home_bias) begin
                    f6_CH_A_d=f6_CH_A_q-home_step;
                end else if (f6_CH_A_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_A_d=f6_CH_A_q+home_step; 
                end 
            end
            2'b01: begin // this is a CHANNEL C
                if (f6_CH_C_q>home_bias) begin
                    f6_CH_C_d=f6_CH_C_q-home_step;
                end else if (f6_CH_C_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_C_d=f6_CH_C_q+home_step;
                end 
            end
            2'b10: begin // this is a CHANNEL B
                if (f6_CH_B_q>home_bias) begin
                    f6_CH_B_d=f6_CH_B_q-home_step;
                end else if (f6_CH_B_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_B_d=f6_CH_B_q+home_step; 
                end 
            end
            2'b11: begin // this is a CHANNEL D
                if (f6_CH_D_q>home_bias) begin
                    f6_CH_D_d=f6_CH_D_q-home_step;
                end else if (f6_CH_D_q<=home_bias) begin //if (CH_A_q<CH_C_q) begin
                    f6_CH_D_d=f6_CH_D_q+home_step; 
                end 
            end
            default: begin
            end
        endcase
    end else begin // if NOT go home
        // F1
        case (f1_addr[2:1])
            2'b00: begin
                f1_CH_A_d= {rom_data[f1_addrs], 8'b10000000};
            end
            2'b01: begin
                f1_CH_C_d= {f1_antidata, 8'b10000000};
            end
            2'b10: begin
                f1_CH_B_d= {rom_data[f1_addrs], 8'b10000000};
            end
            2'b11: begin
                f1_CH_D_d= {f1_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F2
        case (f2_addr[2:1])
            2'b00: begin
                f2_CH_A_d= {rom_data[f2_addrs], 8'b10000000};
            end
            2'b01: begin
                f2_CH_C_d= {f2_antidata, 8'b10000000};
            end
            2'b10: begin
                f2_CH_B_d= {rom_data[f2_addrs],8'b10000000};
            end
            2'b11: begin
                f2_CH_D_d= {f2_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F3
        case (f3_addr[2:1])
            2'b00: begin
                f3_CH_A_d= {rom_data[f3_addrs], 8'b10000000};
            end
            2'b01: begin
                f3_CH_C_d= {f3_antidata, 8'b10000000};
            end
            2'b10: begin
                f3_CH_B_d= {rom_data[f3_addrs], 8'b10000000};
            end
            2'b11: begin
                f3_CH_D_d= {f3_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F4
        case (f4_addr[2:1])
            2'b00: begin
                f4_CH_A_d= {rom_data[f4_addrs],8'b10000000};
            end
            2'b01: begin
                f4_CH_C_d= {f4_antidata, 8'b10000000};
            end
            2'b10: begin
                f4_CH_B_d= {rom_data[f4_addrs],8'b10000000};
            end
            2'b11: begin
                f4_CH_D_d= {f4_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F5
        case (f5_addr[2:1])
            2'b00: begin
                f5_CH_A_d= {rom_data[f5_addrs],8'b10000000};
            end
            2'b01: begin
                f5_CH_C_d= {f5_antidata, 8'b10000000};
            end
            2'b10: begin
                f5_CH_B_d= {rom_data[f5_addrs],8'b10000000};
            end
            2'b11: begin
                f5_CH_D_d= {f5_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase
        // F6
        case (f6_addr[2:1])
            2'b00: begin
                f6_CH_A_d= {rom_data[f6_addrs],8'b10000000};
            end
            2'b01: begin
                f6_CH_C_d= {f6_antidata, 8'b10000000};
            end
            2'b10: begin
                f6_CH_B_d= {rom_data[f6_addrs],8'b10000000};
            end
            2'b11: begin
                f6_CH_D_d= {f6_antidata, 8'b10000000};
            end
        default: begin
            end
        endcase

    end // if go home 

end // always

always @(*) begin
    f1_antidata = 8'hB4 - rom_data[f1_addrs];

    f2_antidata = 8'hB4 - rom_data[f2_addrs];
  f3_antidata = 8'hB4 - rom_data[f3_addrs];
  f4_antidata = 8'hB4 - rom_data[f4_addrs];
  f5_antidata = 8'hB4 - rom_data[f5_addrs];
  f6_antidata = 8'hB4 - rom_data[f6_addrs];

 


  // F1   
  if (f1_addr==0) begin
    f1_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f1_addr==1) begin
    f1_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f1_addr[0]==1'b0) begin
    f1_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f1_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f1_data_d = {6'b000110, f1_addr[2:1], f1_CH_D_q};
            end
            default: begin
            end
        endcase
   end // if addr=0
  // F2
  if (f2_addr==0) begin
    f2_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f2_addr==1) begin
    f2_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f2_addr[0]==1'b0) begin
    f2_data_d = 24'b00111000_0000000000000000; // Vref send in 50% samples  
  end else begin //data in 50%
        case (f2_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f2_data_d = {6'b000110, f2_addr[2:1], f2_CH_D_q};
            end
            default: begin
            end
        endcase
   end // if addr=0
  // F3
  if (f3_addr==0) begin
    f3_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f3_addr==1) begin
    f3_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f3_addr[0]==1'b0) begin
    f3_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f3_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f3_data_d = {6'b000110, f3_addr[2:1], f3_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F4
  if (f4_addr==0) begin
    f4_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f4_addr==1) begin
    f4_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f4_addr[0]==1'b0) begin
    f4_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f4_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f4_data_d = {6'b000110, f4_addr[2:1], f4_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F5
  if (f5_addr==0) begin
    f5_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f5_addr==1) begin
    f5_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f5_addr[0]==1'b0) begin
    f5_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f5_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f5_data_d = {6'b000110, f5_addr[2:1], f5_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
  // F6
  if (f6_addr==0) begin
    f6_data_d = 24'b001010000000000000000001; // set SOFT_RESET once only (in mems cotrol arrd->8)
  end else if (f6_addr==1) begin
    f6_data_d = 24'b00111000_0000000000000000;    // set Vref only once
  end else if (f6_addr[0]==1'b0) begin
    f6_data_d = 24'b00111000_0000000000000000; //Vref send in 50% samples  
  end else begin //data in 50%
        case (f6_addr[2:1])
            2'b00: begin // this is a CHANNEL A
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_A_q};
            end
            2'b01: begin // this is a CHANNEL C
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_C_q};
            end
            2'b10: begin // this is a CHANNEL B
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_B_q};
            end
            2'b11: begin // this is a CHANNEL D
                f6_data_d = {6'b000110, f6_addr[2:1], f6_CH_D_q};
            end
            default: begin
            end
        endcase
  end // if addr=0
end // always

always @(posedge f1_addr[0]) begin
    f1_CH_A_q<=f1_CH_A_d;
    f1_CH_B_q<=f1_CH_B_d;
    f1_CH_C_q<=f1_CH_C_d;
    f1_CH_D_q<=f1_CH_D_d;
end

always @(posedge f2_addr[0]) begin
    f2_CH_A_q<=f2_CH_A_d;
    f2_CH_B_q<=f2_CH_B_d;
    f2_CH_C_q<=f2_CH_C_d;
    f2_CH_D_q<=f2_CH_D_d;
end

always @(posedge f3_addr[0]) begin
    f3_CH_A_q<=f3_CH_A_d;
    f3_CH_B_q<=f3_CH_B_d;
    f3_CH_C_q<=f3_CH_C_d;
    f3_CH_D_q<=f3_CH_D_d;
end

always @(posedge f4_addr[0]) begin
    f4_CH_A_q<=f4_CH_A_d;
    f4_CH_B_q<=f4_CH_B_d;
    f4_CH_C_q<=f4_CH_C_d;
    f4_CH_D_q<=f4_CH_D_d;
end

always @(posedge f5_addr[0]) begin
    f5_CH_A_q<=f5_CH_A_d;
    f5_CH_B_q<=f5_CH_B_d;
    f5_CH_C_q<=f5_CH_C_d;
    f5_CH_D_q<=f5_CH_D_d;
end

always @(posedge f6_addr[0]) begin
    f6_CH_A_q<=f6_CH_A_d;
    f6_CH_B_q<=f6_CH_B_d;
    f6_CH_C_q<=f6_CH_C_d;
    f6_CH_D_q<=f6_CH_D_d;
end

always @(posedge clk) begin
    f1_data_q <= f1_data_d;
    f2_data_q <= f2_data_d;
    f3_data_q <= f3_data_d;
    f4_data_q <= f4_data_d;
    f5_data_q <= f5_data_d;
    f6_data_q <= f6_data_d;
end // always
 
endmodule